magic
tech gf180mcuD
magscale 1 10
timestamp 1755278675
<< mimcap >>
rect -22883 5640 -18883 5720
rect -22883 3800 -22803 5640
rect -18963 3800 -18883 5640
rect -22883 3720 -18883 3800
rect -18269 5640 -14269 5720
rect -18269 3800 -18189 5640
rect -14349 3800 -14269 5640
rect -18269 3720 -14269 3800
rect -13655 5640 -9655 5720
rect -13655 3800 -13575 5640
rect -9735 3800 -9655 5640
rect -13655 3720 -9655 3800
rect -9041 5640 -5041 5720
rect -9041 3800 -8961 5640
rect -5121 3800 -5041 5640
rect -9041 3720 -5041 3800
rect -4427 5640 -427 5720
rect -4427 3800 -4347 5640
rect -507 3800 -427 5640
rect -4427 3720 -427 3800
rect 187 5640 4187 5720
rect 187 3800 267 5640
rect 4107 3800 4187 5640
rect 187 3720 4187 3800
rect 4801 5640 8801 5720
rect 4801 3800 4881 5640
rect 8721 3800 8801 5640
rect 4801 3720 8801 3800
rect 9415 5640 13415 5720
rect 9415 3800 9495 5640
rect 13335 3800 13415 5640
rect 9415 3720 13415 3800
rect 14029 5640 18029 5720
rect 14029 3800 14109 5640
rect 17949 3800 18029 5640
rect 14029 3720 18029 3800
rect 18643 5640 22643 5720
rect 18643 3800 18723 5640
rect 22563 3800 22643 5640
rect 18643 3720 22643 3800
rect -22883 3280 -18883 3360
rect -22883 1440 -22803 3280
rect -18963 1440 -18883 3280
rect -22883 1360 -18883 1440
rect -18269 3280 -14269 3360
rect -18269 1440 -18189 3280
rect -14349 1440 -14269 3280
rect -18269 1360 -14269 1440
rect -13655 3280 -9655 3360
rect -13655 1440 -13575 3280
rect -9735 1440 -9655 3280
rect -13655 1360 -9655 1440
rect -9041 3280 -5041 3360
rect -9041 1440 -8961 3280
rect -5121 1440 -5041 3280
rect -9041 1360 -5041 1440
rect -4427 3280 -427 3360
rect -4427 1440 -4347 3280
rect -507 1440 -427 3280
rect -4427 1360 -427 1440
rect 187 3280 4187 3360
rect 187 1440 267 3280
rect 4107 1440 4187 3280
rect 187 1360 4187 1440
rect 4801 3280 8801 3360
rect 4801 1440 4881 3280
rect 8721 1440 8801 3280
rect 4801 1360 8801 1440
rect 9415 3280 13415 3360
rect 9415 1440 9495 3280
rect 13335 1440 13415 3280
rect 9415 1360 13415 1440
rect 14029 3280 18029 3360
rect 14029 1440 14109 3280
rect 17949 1440 18029 3280
rect 14029 1360 18029 1440
rect 18643 3280 22643 3360
rect 18643 1440 18723 3280
rect 22563 1440 22643 3280
rect 18643 1360 22643 1440
rect -22883 920 -18883 1000
rect -22883 -920 -22803 920
rect -18963 -920 -18883 920
rect -22883 -1000 -18883 -920
rect -18269 920 -14269 1000
rect -18269 -920 -18189 920
rect -14349 -920 -14269 920
rect -18269 -1000 -14269 -920
rect -13655 920 -9655 1000
rect -13655 -920 -13575 920
rect -9735 -920 -9655 920
rect -13655 -1000 -9655 -920
rect -9041 920 -5041 1000
rect -9041 -920 -8961 920
rect -5121 -920 -5041 920
rect -9041 -1000 -5041 -920
rect -4427 920 -427 1000
rect -4427 -920 -4347 920
rect -507 -920 -427 920
rect -4427 -1000 -427 -920
rect 187 920 4187 1000
rect 187 -920 267 920
rect 4107 -920 4187 920
rect 187 -1000 4187 -920
rect 4801 920 8801 1000
rect 4801 -920 4881 920
rect 8721 -920 8801 920
rect 4801 -1000 8801 -920
rect 9415 920 13415 1000
rect 9415 -920 9495 920
rect 13335 -920 13415 920
rect 9415 -1000 13415 -920
rect 14029 920 18029 1000
rect 14029 -920 14109 920
rect 17949 -920 18029 920
rect 14029 -1000 18029 -920
rect 18643 920 22643 1000
rect 18643 -920 18723 920
rect 22563 -920 22643 920
rect 18643 -1000 22643 -920
rect -22883 -1440 -18883 -1360
rect -22883 -3280 -22803 -1440
rect -18963 -3280 -18883 -1440
rect -22883 -3360 -18883 -3280
rect -18269 -1440 -14269 -1360
rect -18269 -3280 -18189 -1440
rect -14349 -3280 -14269 -1440
rect -18269 -3360 -14269 -3280
rect -13655 -1440 -9655 -1360
rect -13655 -3280 -13575 -1440
rect -9735 -3280 -9655 -1440
rect -13655 -3360 -9655 -3280
rect -9041 -1440 -5041 -1360
rect -9041 -3280 -8961 -1440
rect -5121 -3280 -5041 -1440
rect -9041 -3360 -5041 -3280
rect -4427 -1440 -427 -1360
rect -4427 -3280 -4347 -1440
rect -507 -3280 -427 -1440
rect -4427 -3360 -427 -3280
rect 187 -1440 4187 -1360
rect 187 -3280 267 -1440
rect 4107 -3280 4187 -1440
rect 187 -3360 4187 -3280
rect 4801 -1440 8801 -1360
rect 4801 -3280 4881 -1440
rect 8721 -3280 8801 -1440
rect 4801 -3360 8801 -3280
rect 9415 -1440 13415 -1360
rect 9415 -3280 9495 -1440
rect 13335 -3280 13415 -1440
rect 9415 -3360 13415 -3280
rect 14029 -1440 18029 -1360
rect 14029 -3280 14109 -1440
rect 17949 -3280 18029 -1440
rect 14029 -3360 18029 -3280
rect 18643 -1440 22643 -1360
rect 18643 -3280 18723 -1440
rect 22563 -3280 22643 -1440
rect 18643 -3360 22643 -3280
rect -22883 -3800 -18883 -3720
rect -22883 -5640 -22803 -3800
rect -18963 -5640 -18883 -3800
rect -22883 -5720 -18883 -5640
rect -18269 -3800 -14269 -3720
rect -18269 -5640 -18189 -3800
rect -14349 -5640 -14269 -3800
rect -18269 -5720 -14269 -5640
rect -13655 -3800 -9655 -3720
rect -13655 -5640 -13575 -3800
rect -9735 -5640 -9655 -3800
rect -13655 -5720 -9655 -5640
rect -9041 -3800 -5041 -3720
rect -9041 -5640 -8961 -3800
rect -5121 -5640 -5041 -3800
rect -9041 -5720 -5041 -5640
rect -4427 -3800 -427 -3720
rect -4427 -5640 -4347 -3800
rect -507 -5640 -427 -3800
rect -4427 -5720 -427 -5640
rect 187 -3800 4187 -3720
rect 187 -5640 267 -3800
rect 4107 -5640 4187 -3800
rect 187 -5720 4187 -5640
rect 4801 -3800 8801 -3720
rect 4801 -5640 4881 -3800
rect 8721 -5640 8801 -3800
rect 4801 -5720 8801 -5640
rect 9415 -3800 13415 -3720
rect 9415 -5640 9495 -3800
rect 13335 -5640 13415 -3800
rect 9415 -5720 13415 -5640
rect 14029 -3800 18029 -3720
rect 14029 -5640 14109 -3800
rect 17949 -5640 18029 -3800
rect 14029 -5720 18029 -5640
rect 18643 -3800 22643 -3720
rect 18643 -5640 18723 -3800
rect 22563 -5640 22643 -3800
rect 18643 -5720 22643 -5640
<< mimcapcontact >>
rect -22803 3800 -18963 5640
rect -18189 3800 -14349 5640
rect -13575 3800 -9735 5640
rect -8961 3800 -5121 5640
rect -4347 3800 -507 5640
rect 267 3800 4107 5640
rect 4881 3800 8721 5640
rect 9495 3800 13335 5640
rect 14109 3800 17949 5640
rect 18723 3800 22563 5640
rect -22803 1440 -18963 3280
rect -18189 1440 -14349 3280
rect -13575 1440 -9735 3280
rect -8961 1440 -5121 3280
rect -4347 1440 -507 3280
rect 267 1440 4107 3280
rect 4881 1440 8721 3280
rect 9495 1440 13335 3280
rect 14109 1440 17949 3280
rect 18723 1440 22563 3280
rect -22803 -920 -18963 920
rect -18189 -920 -14349 920
rect -13575 -920 -9735 920
rect -8961 -920 -5121 920
rect -4347 -920 -507 920
rect 267 -920 4107 920
rect 4881 -920 8721 920
rect 9495 -920 13335 920
rect 14109 -920 17949 920
rect 18723 -920 22563 920
rect -22803 -3280 -18963 -1440
rect -18189 -3280 -14349 -1440
rect -13575 -3280 -9735 -1440
rect -8961 -3280 -5121 -1440
rect -4347 -3280 -507 -1440
rect 267 -3280 4107 -1440
rect 4881 -3280 8721 -1440
rect 9495 -3280 13335 -1440
rect 14109 -3280 17949 -1440
rect 18723 -3280 22563 -1440
rect -22803 -5640 -18963 -3800
rect -18189 -5640 -14349 -3800
rect -13575 -5640 -9735 -3800
rect -8961 -5640 -5121 -3800
rect -4347 -5640 -507 -3800
rect 267 -5640 4107 -3800
rect 4881 -5640 8721 -3800
rect 9495 -5640 13335 -3800
rect 14109 -5640 17949 -3800
rect 18723 -5640 22563 -3800
<< metal4 >>
rect -23003 5773 -18523 5840
rect -23003 5720 -18673 5773
rect -23003 3720 -22883 5720
rect -18883 3720 -18673 5720
rect -23003 3667 -18673 3720
rect -18585 3667 -18523 5773
rect -23003 3600 -18523 3667
rect -18389 5773 -13909 5840
rect -18389 5720 -14059 5773
rect -18389 3720 -18269 5720
rect -14269 3720 -14059 5720
rect -18389 3667 -14059 3720
rect -13971 3667 -13909 5773
rect -18389 3600 -13909 3667
rect -13775 5773 -9295 5840
rect -13775 5720 -9445 5773
rect -13775 3720 -13655 5720
rect -9655 3720 -9445 5720
rect -13775 3667 -9445 3720
rect -9357 3667 -9295 5773
rect -13775 3600 -9295 3667
rect -9161 5773 -4681 5840
rect -9161 5720 -4831 5773
rect -9161 3720 -9041 5720
rect -5041 3720 -4831 5720
rect -9161 3667 -4831 3720
rect -4743 3667 -4681 5773
rect -9161 3600 -4681 3667
rect -4547 5773 -67 5840
rect -4547 5720 -217 5773
rect -4547 3720 -4427 5720
rect -427 3720 -217 5720
rect -4547 3667 -217 3720
rect -129 3667 -67 5773
rect -4547 3600 -67 3667
rect 67 5773 4547 5840
rect 67 5720 4397 5773
rect 67 3720 187 5720
rect 4187 3720 4397 5720
rect 67 3667 4397 3720
rect 4485 3667 4547 5773
rect 67 3600 4547 3667
rect 4681 5773 9161 5840
rect 4681 5720 9011 5773
rect 4681 3720 4801 5720
rect 8801 3720 9011 5720
rect 4681 3667 9011 3720
rect 9099 3667 9161 5773
rect 4681 3600 9161 3667
rect 9295 5773 13775 5840
rect 9295 5720 13625 5773
rect 9295 3720 9415 5720
rect 13415 3720 13625 5720
rect 9295 3667 13625 3720
rect 13713 3667 13775 5773
rect 9295 3600 13775 3667
rect 13909 5773 18389 5840
rect 13909 5720 18239 5773
rect 13909 3720 14029 5720
rect 18029 3720 18239 5720
rect 13909 3667 18239 3720
rect 18327 3667 18389 5773
rect 13909 3600 18389 3667
rect 18523 5773 23003 5840
rect 18523 5720 22853 5773
rect 18523 3720 18643 5720
rect 22643 3720 22853 5720
rect 18523 3667 22853 3720
rect 22941 3667 23003 5773
rect 18523 3600 23003 3667
rect -23003 3413 -18523 3480
rect -23003 3360 -18673 3413
rect -23003 1360 -22883 3360
rect -18883 1360 -18673 3360
rect -23003 1307 -18673 1360
rect -18585 1307 -18523 3413
rect -23003 1240 -18523 1307
rect -18389 3413 -13909 3480
rect -18389 3360 -14059 3413
rect -18389 1360 -18269 3360
rect -14269 1360 -14059 3360
rect -18389 1307 -14059 1360
rect -13971 1307 -13909 3413
rect -18389 1240 -13909 1307
rect -13775 3413 -9295 3480
rect -13775 3360 -9445 3413
rect -13775 1360 -13655 3360
rect -9655 1360 -9445 3360
rect -13775 1307 -9445 1360
rect -9357 1307 -9295 3413
rect -13775 1240 -9295 1307
rect -9161 3413 -4681 3480
rect -9161 3360 -4831 3413
rect -9161 1360 -9041 3360
rect -5041 1360 -4831 3360
rect -9161 1307 -4831 1360
rect -4743 1307 -4681 3413
rect -9161 1240 -4681 1307
rect -4547 3413 -67 3480
rect -4547 3360 -217 3413
rect -4547 1360 -4427 3360
rect -427 1360 -217 3360
rect -4547 1307 -217 1360
rect -129 1307 -67 3413
rect -4547 1240 -67 1307
rect 67 3413 4547 3480
rect 67 3360 4397 3413
rect 67 1360 187 3360
rect 4187 1360 4397 3360
rect 67 1307 4397 1360
rect 4485 1307 4547 3413
rect 67 1240 4547 1307
rect 4681 3413 9161 3480
rect 4681 3360 9011 3413
rect 4681 1360 4801 3360
rect 8801 1360 9011 3360
rect 4681 1307 9011 1360
rect 9099 1307 9161 3413
rect 4681 1240 9161 1307
rect 9295 3413 13775 3480
rect 9295 3360 13625 3413
rect 9295 1360 9415 3360
rect 13415 1360 13625 3360
rect 9295 1307 13625 1360
rect 13713 1307 13775 3413
rect 9295 1240 13775 1307
rect 13909 3413 18389 3480
rect 13909 3360 18239 3413
rect 13909 1360 14029 3360
rect 18029 1360 18239 3360
rect 13909 1307 18239 1360
rect 18327 1307 18389 3413
rect 13909 1240 18389 1307
rect 18523 3413 23003 3480
rect 18523 3360 22853 3413
rect 18523 1360 18643 3360
rect 22643 1360 22853 3360
rect 18523 1307 22853 1360
rect 22941 1307 23003 3413
rect 18523 1240 23003 1307
rect -23003 1053 -18523 1120
rect -23003 1000 -18673 1053
rect -23003 -1000 -22883 1000
rect -18883 -1000 -18673 1000
rect -23003 -1053 -18673 -1000
rect -18585 -1053 -18523 1053
rect -23003 -1120 -18523 -1053
rect -18389 1053 -13909 1120
rect -18389 1000 -14059 1053
rect -18389 -1000 -18269 1000
rect -14269 -1000 -14059 1000
rect -18389 -1053 -14059 -1000
rect -13971 -1053 -13909 1053
rect -18389 -1120 -13909 -1053
rect -13775 1053 -9295 1120
rect -13775 1000 -9445 1053
rect -13775 -1000 -13655 1000
rect -9655 -1000 -9445 1000
rect -13775 -1053 -9445 -1000
rect -9357 -1053 -9295 1053
rect -13775 -1120 -9295 -1053
rect -9161 1053 -4681 1120
rect -9161 1000 -4831 1053
rect -9161 -1000 -9041 1000
rect -5041 -1000 -4831 1000
rect -9161 -1053 -4831 -1000
rect -4743 -1053 -4681 1053
rect -9161 -1120 -4681 -1053
rect -4547 1053 -67 1120
rect -4547 1000 -217 1053
rect -4547 -1000 -4427 1000
rect -427 -1000 -217 1000
rect -4547 -1053 -217 -1000
rect -129 -1053 -67 1053
rect -4547 -1120 -67 -1053
rect 67 1053 4547 1120
rect 67 1000 4397 1053
rect 67 -1000 187 1000
rect 4187 -1000 4397 1000
rect 67 -1053 4397 -1000
rect 4485 -1053 4547 1053
rect 67 -1120 4547 -1053
rect 4681 1053 9161 1120
rect 4681 1000 9011 1053
rect 4681 -1000 4801 1000
rect 8801 -1000 9011 1000
rect 4681 -1053 9011 -1000
rect 9099 -1053 9161 1053
rect 4681 -1120 9161 -1053
rect 9295 1053 13775 1120
rect 9295 1000 13625 1053
rect 9295 -1000 9415 1000
rect 13415 -1000 13625 1000
rect 9295 -1053 13625 -1000
rect 13713 -1053 13775 1053
rect 9295 -1120 13775 -1053
rect 13909 1053 18389 1120
rect 13909 1000 18239 1053
rect 13909 -1000 14029 1000
rect 18029 -1000 18239 1000
rect 13909 -1053 18239 -1000
rect 18327 -1053 18389 1053
rect 13909 -1120 18389 -1053
rect 18523 1053 23003 1120
rect 18523 1000 22853 1053
rect 18523 -1000 18643 1000
rect 22643 -1000 22853 1000
rect 18523 -1053 22853 -1000
rect 22941 -1053 23003 1053
rect 18523 -1120 23003 -1053
rect -23003 -1307 -18523 -1240
rect -23003 -1360 -18673 -1307
rect -23003 -3360 -22883 -1360
rect -18883 -3360 -18673 -1360
rect -23003 -3413 -18673 -3360
rect -18585 -3413 -18523 -1307
rect -23003 -3480 -18523 -3413
rect -18389 -1307 -13909 -1240
rect -18389 -1360 -14059 -1307
rect -18389 -3360 -18269 -1360
rect -14269 -3360 -14059 -1360
rect -18389 -3413 -14059 -3360
rect -13971 -3413 -13909 -1307
rect -18389 -3480 -13909 -3413
rect -13775 -1307 -9295 -1240
rect -13775 -1360 -9445 -1307
rect -13775 -3360 -13655 -1360
rect -9655 -3360 -9445 -1360
rect -13775 -3413 -9445 -3360
rect -9357 -3413 -9295 -1307
rect -13775 -3480 -9295 -3413
rect -9161 -1307 -4681 -1240
rect -9161 -1360 -4831 -1307
rect -9161 -3360 -9041 -1360
rect -5041 -3360 -4831 -1360
rect -9161 -3413 -4831 -3360
rect -4743 -3413 -4681 -1307
rect -9161 -3480 -4681 -3413
rect -4547 -1307 -67 -1240
rect -4547 -1360 -217 -1307
rect -4547 -3360 -4427 -1360
rect -427 -3360 -217 -1360
rect -4547 -3413 -217 -3360
rect -129 -3413 -67 -1307
rect -4547 -3480 -67 -3413
rect 67 -1307 4547 -1240
rect 67 -1360 4397 -1307
rect 67 -3360 187 -1360
rect 4187 -3360 4397 -1360
rect 67 -3413 4397 -3360
rect 4485 -3413 4547 -1307
rect 67 -3480 4547 -3413
rect 4681 -1307 9161 -1240
rect 4681 -1360 9011 -1307
rect 4681 -3360 4801 -1360
rect 8801 -3360 9011 -1360
rect 4681 -3413 9011 -3360
rect 9099 -3413 9161 -1307
rect 4681 -3480 9161 -3413
rect 9295 -1307 13775 -1240
rect 9295 -1360 13625 -1307
rect 9295 -3360 9415 -1360
rect 13415 -3360 13625 -1360
rect 9295 -3413 13625 -3360
rect 13713 -3413 13775 -1307
rect 9295 -3480 13775 -3413
rect 13909 -1307 18389 -1240
rect 13909 -1360 18239 -1307
rect 13909 -3360 14029 -1360
rect 18029 -3360 18239 -1360
rect 13909 -3413 18239 -3360
rect 18327 -3413 18389 -1307
rect 13909 -3480 18389 -3413
rect 18523 -1307 23003 -1240
rect 18523 -1360 22853 -1307
rect 18523 -3360 18643 -1360
rect 22643 -3360 22853 -1360
rect 18523 -3413 22853 -3360
rect 22941 -3413 23003 -1307
rect 18523 -3480 23003 -3413
rect -23003 -3667 -18523 -3600
rect -23003 -3720 -18673 -3667
rect -23003 -5720 -22883 -3720
rect -18883 -5720 -18673 -3720
rect -23003 -5773 -18673 -5720
rect -18585 -5773 -18523 -3667
rect -23003 -5840 -18523 -5773
rect -18389 -3667 -13909 -3600
rect -18389 -3720 -14059 -3667
rect -18389 -5720 -18269 -3720
rect -14269 -5720 -14059 -3720
rect -18389 -5773 -14059 -5720
rect -13971 -5773 -13909 -3667
rect -18389 -5840 -13909 -5773
rect -13775 -3667 -9295 -3600
rect -13775 -3720 -9445 -3667
rect -13775 -5720 -13655 -3720
rect -9655 -5720 -9445 -3720
rect -13775 -5773 -9445 -5720
rect -9357 -5773 -9295 -3667
rect -13775 -5840 -9295 -5773
rect -9161 -3667 -4681 -3600
rect -9161 -3720 -4831 -3667
rect -9161 -5720 -9041 -3720
rect -5041 -5720 -4831 -3720
rect -9161 -5773 -4831 -5720
rect -4743 -5773 -4681 -3667
rect -9161 -5840 -4681 -5773
rect -4547 -3667 -67 -3600
rect -4547 -3720 -217 -3667
rect -4547 -5720 -4427 -3720
rect -427 -5720 -217 -3720
rect -4547 -5773 -217 -5720
rect -129 -5773 -67 -3667
rect -4547 -5840 -67 -5773
rect 67 -3667 4547 -3600
rect 67 -3720 4397 -3667
rect 67 -5720 187 -3720
rect 4187 -5720 4397 -3720
rect 67 -5773 4397 -5720
rect 4485 -5773 4547 -3667
rect 67 -5840 4547 -5773
rect 4681 -3667 9161 -3600
rect 4681 -3720 9011 -3667
rect 4681 -5720 4801 -3720
rect 8801 -5720 9011 -3720
rect 4681 -5773 9011 -5720
rect 9099 -5773 9161 -3667
rect 4681 -5840 9161 -5773
rect 9295 -3667 13775 -3600
rect 9295 -3720 13625 -3667
rect 9295 -5720 9415 -3720
rect 13415 -5720 13625 -3720
rect 9295 -5773 13625 -5720
rect 13713 -5773 13775 -3667
rect 9295 -5840 13775 -5773
rect 13909 -3667 18389 -3600
rect 13909 -3720 18239 -3667
rect 13909 -5720 14029 -3720
rect 18029 -5720 18239 -3720
rect 13909 -5773 18239 -5720
rect 18327 -5773 18389 -3667
rect 13909 -5840 18389 -5773
rect 18523 -3667 23003 -3600
rect 18523 -3720 22853 -3667
rect 18523 -5720 18643 -3720
rect 22643 -5720 22853 -3720
rect 18523 -5773 22853 -5720
rect 22941 -5773 23003 -3667
rect 18523 -5840 23003 -5773
<< via4 >>
rect -18673 3667 -18585 5773
rect -14059 3667 -13971 5773
rect -9445 3667 -9357 5773
rect -4831 3667 -4743 5773
rect -217 3667 -129 5773
rect 4397 3667 4485 5773
rect 9011 3667 9099 5773
rect 13625 3667 13713 5773
rect 18239 3667 18327 5773
rect 22853 3667 22941 5773
rect -18673 1307 -18585 3413
rect -14059 1307 -13971 3413
rect -9445 1307 -9357 3413
rect -4831 1307 -4743 3413
rect -217 1307 -129 3413
rect 4397 1307 4485 3413
rect 9011 1307 9099 3413
rect 13625 1307 13713 3413
rect 18239 1307 18327 3413
rect 22853 1307 22941 3413
rect -18673 -1053 -18585 1053
rect -14059 -1053 -13971 1053
rect -9445 -1053 -9357 1053
rect -4831 -1053 -4743 1053
rect -217 -1053 -129 1053
rect 4397 -1053 4485 1053
rect 9011 -1053 9099 1053
rect 13625 -1053 13713 1053
rect 18239 -1053 18327 1053
rect 22853 -1053 22941 1053
rect -18673 -3413 -18585 -1307
rect -14059 -3413 -13971 -1307
rect -9445 -3413 -9357 -1307
rect -4831 -3413 -4743 -1307
rect -217 -3413 -129 -1307
rect 4397 -3413 4485 -1307
rect 9011 -3413 9099 -1307
rect 13625 -3413 13713 -1307
rect 18239 -3413 18327 -1307
rect 22853 -3413 22941 -1307
rect -18673 -5773 -18585 -3667
rect -14059 -5773 -13971 -3667
rect -9445 -5773 -9357 -3667
rect -4831 -5773 -4743 -3667
rect -217 -5773 -129 -3667
rect 4397 -5773 4485 -3667
rect 9011 -5773 9099 -3667
rect 13625 -5773 13713 -3667
rect 18239 -5773 18327 -3667
rect 22853 -5773 22941 -3667
<< metal5 >>
rect -20989 5640 -20777 5900
rect -18735 5773 -18523 5900
rect -20989 3280 -20777 3800
rect -18735 3667 -18673 5773
rect -18585 3667 -18523 5773
rect -16375 5640 -16163 5900
rect -14121 5773 -13909 5900
rect -18735 3413 -18523 3667
rect -20989 920 -20777 1440
rect -18735 1307 -18673 3413
rect -18585 1307 -18523 3413
rect -16375 3280 -16163 3800
rect -14121 3667 -14059 5773
rect -13971 3667 -13909 5773
rect -11761 5640 -11549 5900
rect -9507 5773 -9295 5900
rect -14121 3413 -13909 3667
rect -18735 1053 -18523 1307
rect -20989 -1440 -20777 -920
rect -18735 -1053 -18673 1053
rect -18585 -1053 -18523 1053
rect -16375 920 -16163 1440
rect -14121 1307 -14059 3413
rect -13971 1307 -13909 3413
rect -11761 3280 -11549 3800
rect -9507 3667 -9445 5773
rect -9357 3667 -9295 5773
rect -7147 5640 -6935 5900
rect -4893 5773 -4681 5900
rect -9507 3413 -9295 3667
rect -14121 1053 -13909 1307
rect -18735 -1307 -18523 -1053
rect -20989 -3800 -20777 -3280
rect -18735 -3413 -18673 -1307
rect -18585 -3413 -18523 -1307
rect -16375 -1440 -16163 -920
rect -14121 -1053 -14059 1053
rect -13971 -1053 -13909 1053
rect -11761 920 -11549 1440
rect -9507 1307 -9445 3413
rect -9357 1307 -9295 3413
rect -7147 3280 -6935 3800
rect -4893 3667 -4831 5773
rect -4743 3667 -4681 5773
rect -2533 5640 -2321 5900
rect -279 5773 -67 5900
rect -4893 3413 -4681 3667
rect -9507 1053 -9295 1307
rect -14121 -1307 -13909 -1053
rect -18735 -3667 -18523 -3413
rect -20989 -5900 -20777 -5640
rect -18735 -5773 -18673 -3667
rect -18585 -5773 -18523 -3667
rect -16375 -3800 -16163 -3280
rect -14121 -3413 -14059 -1307
rect -13971 -3413 -13909 -1307
rect -11761 -1440 -11549 -920
rect -9507 -1053 -9445 1053
rect -9357 -1053 -9295 1053
rect -7147 920 -6935 1440
rect -4893 1307 -4831 3413
rect -4743 1307 -4681 3413
rect -2533 3280 -2321 3800
rect -279 3667 -217 5773
rect -129 3667 -67 5773
rect 2081 5640 2293 5900
rect 4335 5773 4547 5900
rect -279 3413 -67 3667
rect -4893 1053 -4681 1307
rect -9507 -1307 -9295 -1053
rect -14121 -3667 -13909 -3413
rect -18735 -5900 -18523 -5773
rect -16375 -5900 -16163 -5640
rect -14121 -5773 -14059 -3667
rect -13971 -5773 -13909 -3667
rect -11761 -3800 -11549 -3280
rect -9507 -3413 -9445 -1307
rect -9357 -3413 -9295 -1307
rect -7147 -1440 -6935 -920
rect -4893 -1053 -4831 1053
rect -4743 -1053 -4681 1053
rect -2533 920 -2321 1440
rect -279 1307 -217 3413
rect -129 1307 -67 3413
rect 2081 3280 2293 3800
rect 4335 3667 4397 5773
rect 4485 3667 4547 5773
rect 6695 5640 6907 5900
rect 8949 5773 9161 5900
rect 4335 3413 4547 3667
rect -279 1053 -67 1307
rect -4893 -1307 -4681 -1053
rect -9507 -3667 -9295 -3413
rect -14121 -5900 -13909 -5773
rect -11761 -5900 -11549 -5640
rect -9507 -5773 -9445 -3667
rect -9357 -5773 -9295 -3667
rect -7147 -3800 -6935 -3280
rect -4893 -3413 -4831 -1307
rect -4743 -3413 -4681 -1307
rect -2533 -1440 -2321 -920
rect -279 -1053 -217 1053
rect -129 -1053 -67 1053
rect 2081 920 2293 1440
rect 4335 1307 4397 3413
rect 4485 1307 4547 3413
rect 6695 3280 6907 3800
rect 8949 3667 9011 5773
rect 9099 3667 9161 5773
rect 11309 5640 11521 5900
rect 13563 5773 13775 5900
rect 8949 3413 9161 3667
rect 4335 1053 4547 1307
rect -279 -1307 -67 -1053
rect -4893 -3667 -4681 -3413
rect -9507 -5900 -9295 -5773
rect -7147 -5900 -6935 -5640
rect -4893 -5773 -4831 -3667
rect -4743 -5773 -4681 -3667
rect -2533 -3800 -2321 -3280
rect -279 -3413 -217 -1307
rect -129 -3413 -67 -1307
rect 2081 -1440 2293 -920
rect 4335 -1053 4397 1053
rect 4485 -1053 4547 1053
rect 6695 920 6907 1440
rect 8949 1307 9011 3413
rect 9099 1307 9161 3413
rect 11309 3280 11521 3800
rect 13563 3667 13625 5773
rect 13713 3667 13775 5773
rect 15923 5640 16135 5900
rect 18177 5773 18389 5900
rect 13563 3413 13775 3667
rect 8949 1053 9161 1307
rect 4335 -1307 4547 -1053
rect -279 -3667 -67 -3413
rect -4893 -5900 -4681 -5773
rect -2533 -5900 -2321 -5640
rect -279 -5773 -217 -3667
rect -129 -5773 -67 -3667
rect 2081 -3800 2293 -3280
rect 4335 -3413 4397 -1307
rect 4485 -3413 4547 -1307
rect 6695 -1440 6907 -920
rect 8949 -1053 9011 1053
rect 9099 -1053 9161 1053
rect 11309 920 11521 1440
rect 13563 1307 13625 3413
rect 13713 1307 13775 3413
rect 15923 3280 16135 3800
rect 18177 3667 18239 5773
rect 18327 3667 18389 5773
rect 20537 5640 20749 5900
rect 22791 5773 23003 5900
rect 18177 3413 18389 3667
rect 13563 1053 13775 1307
rect 8949 -1307 9161 -1053
rect 4335 -3667 4547 -3413
rect -279 -5900 -67 -5773
rect 2081 -5900 2293 -5640
rect 4335 -5773 4397 -3667
rect 4485 -5773 4547 -3667
rect 6695 -3800 6907 -3280
rect 8949 -3413 9011 -1307
rect 9099 -3413 9161 -1307
rect 11309 -1440 11521 -920
rect 13563 -1053 13625 1053
rect 13713 -1053 13775 1053
rect 15923 920 16135 1440
rect 18177 1307 18239 3413
rect 18327 1307 18389 3413
rect 20537 3280 20749 3800
rect 22791 3667 22853 5773
rect 22941 3667 23003 5773
rect 22791 3413 23003 3667
rect 18177 1053 18389 1307
rect 13563 -1307 13775 -1053
rect 8949 -3667 9161 -3413
rect 4335 -5900 4547 -5773
rect 6695 -5900 6907 -5640
rect 8949 -5773 9011 -3667
rect 9099 -5773 9161 -3667
rect 11309 -3800 11521 -3280
rect 13563 -3413 13625 -1307
rect 13713 -3413 13775 -1307
rect 15923 -1440 16135 -920
rect 18177 -1053 18239 1053
rect 18327 -1053 18389 1053
rect 20537 920 20749 1440
rect 22791 1307 22853 3413
rect 22941 1307 23003 3413
rect 22791 1053 23003 1307
rect 18177 -1307 18389 -1053
rect 13563 -3667 13775 -3413
rect 8949 -5900 9161 -5773
rect 11309 -5900 11521 -5640
rect 13563 -5773 13625 -3667
rect 13713 -5773 13775 -3667
rect 15923 -3800 16135 -3280
rect 18177 -3413 18239 -1307
rect 18327 -3413 18389 -1307
rect 20537 -1440 20749 -920
rect 22791 -1053 22853 1053
rect 22941 -1053 23003 1053
rect 22791 -1307 23003 -1053
rect 18177 -3667 18389 -3413
rect 13563 -5900 13775 -5773
rect 15923 -5900 16135 -5640
rect 18177 -5773 18239 -3667
rect 18327 -5773 18389 -3667
rect 20537 -3800 20749 -3280
rect 22791 -3413 22853 -1307
rect 22941 -3413 23003 -1307
rect 22791 -3667 23003 -3413
rect 18177 -5900 18389 -5773
rect 20537 -5900 20749 -5640
rect 22791 -5773 22853 -3667
rect 22941 -5773 23003 -3667
rect 22791 -5900 23003 -5773
<< properties >>
string FIXED_BBOX 18523 3600 22763 5840
string gencell cap_mim_2p0fF
string library gf180mcu
string parameters w 20 l 10 val 6.2k carea 25.00 cperi 20.00 class capacitor nx 10 ny 5 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 1 tconnect 1
<< end >>
