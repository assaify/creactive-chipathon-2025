* Extracted by KLayout with GF180MCU LVS runset on : 08/09/2025 13:33

.SUBCKT tail_current_diff_out VSS I3C I2C IBIAS I3A I2A I1A I1C I3B I1B I2B
M$1 VSS VSS VSS VSS nfet_03v3 L=0.8U W=75U AS=36.3P AD=36.3P PS=124.36U
+ PD=124.36U
M$2 I2C IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$4 I3C IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$28 I2A IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$30 I3A IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$38 I1A IBIAS VSS VSS nfet_03v3 L=0.8U W=7.5U AS=3P AD=3P PS=9.1U PD=9.1U
M$39 I1A I1A I1A VSS nfet_03v3 L=0.8U W=7.5U AS=3.7875P AD=3.7875P PS=13.27U
+ PD=13.27U
M$40 I1C I1C I1C VSS nfet_03v3 L=0.8U W=7.5U AS=3.7875P AD=3.7875P PS=13.27U
+ PD=13.27U
M$41 VSS IBIAS I1C VSS nfet_03v3 L=0.8U W=7.5U AS=3P AD=3P PS=9.1U PD=9.1U
M$54 I2B IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$56 I3B IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$64 I1B IBIAS VSS VSS nfet_03v3 L=0.8U W=7.5U AS=3P AD=3P PS=9.1U PD=9.1U
M$65 I1B I1B I1B VSS nfet_03v3 L=0.8U W=7.5U AS=3.7875P AD=3.7875P PS=13.27U
+ PD=13.27U
M$66 IBIAS IBIAS IBIAS VSS nfet_03v3 L=0.8U W=7.5U AS=3.7875P AD=3.7875P
+ PS=13.27U PD=13.27U
M$67 VSS IBIAS IBIAS VSS nfet_03v3 L=0.8U W=7.5U AS=3P AD=3P PS=9.1U PD=9.1U
.ENDS tail_current_diff_out
