magic
tech gf180mcuD
magscale 1 10
timestamp 1755276408
<< pwell >>
rect -336 -1308 336 1308
<< psubdiff >>
rect -312 1212 312 1284
rect -312 1168 -240 1212
rect -312 -1168 -299 1168
rect -253 -1168 -240 1168
rect 240 1168 312 1212
rect -312 -1212 -240 -1168
rect 240 -1168 253 1168
rect 299 -1168 312 1168
rect 240 -1212 312 -1168
rect -312 -1284 312 -1212
<< psubdiffcont >>
rect -299 -1168 -253 1168
rect 253 -1168 299 1168
<< polysilicon >>
rect -100 1059 100 1072
rect -100 1013 -87 1059
rect 87 1013 100 1059
rect -100 950 100 1013
rect -100 -1013 100 -950
rect -100 -1059 -87 -1013
rect 87 -1059 100 -1013
rect -100 -1072 100 -1059
<< polycontact >>
rect -87 1013 87 1059
rect -87 -1059 87 -1013
<< nhighres >>
rect -100 -950 100 950
<< metal1 >>
rect -299 1225 299 1271
rect -299 1168 -253 1225
rect 253 1168 299 1225
rect -98 1013 -87 1059
rect 87 1013 98 1059
rect -98 -1059 -87 -1013
rect 87 -1059 98 -1013
rect -299 -1225 -253 -1168
rect 253 -1225 299 -1168
rect -299 -1271 299 -1225
<< properties >>
string FIXED_BBOX -276 -1248 276 1248
string gencell ppolyf_u_1k
string library gf180mcu
string parameters w 1.0 l 9.5 m 1 nx 1 wmin 1.000 lmin 1.000 class resistor rho 1000 val 9.5k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
