magic
tech gf180mcuD
magscale 1 10
timestamp 1758729012
<< error_s >>
rect 6609 31130 6610 31251
rect 11913 31130 11914 31251
rect 6609 28478 6610 28599
rect 11913 28478 11914 28599
rect 6609 25826 6610 25947
rect 11913 25826 11914 25947
rect 6609 23174 6610 23295
rect 11913 23174 11914 23295
rect 6609 20522 6610 20643
rect 11913 20522 11914 20643
rect 6609 17870 6610 17991
rect 11913 17870 11914 17991
rect 6609 15218 6610 15339
rect 11913 15218 11914 15339
rect 6609 12566 6610 12687
rect 11913 12566 11914 12687
rect 6609 9914 6610 10035
rect 11913 9914 11914 10035
rect 6609 7262 6610 7383
rect 11913 7262 11914 7383
rect 6609 4610 6610 4731
rect 11913 4610 11914 4731
<< metal4 >>
rect 4078 34512 4490 35088
rect 6730 34512 7142 35088
rect 9382 34512 9794 35088
rect 12034 34512 12446 35088
rect 576 34496 15948 34512
rect 576 34440 4100 34496
rect 4468 34440 6752 34496
rect 7120 34440 9404 34496
rect 9772 34440 12056 34496
rect 12424 34440 15948 34496
rect 576 34424 15948 34440
rect 576 31010 664 34424
rect 4078 33848 4490 34424
rect 6730 33848 7142 34424
rect 9382 33848 9794 34424
rect 12034 33848 12446 34424
rect 1838 33530 4078 33608
rect 1838 33474 2202 33530
rect 4026 33474 4078 33530
rect 1838 33250 4078 33474
rect 7142 33530 9382 33608
rect 7142 33474 7194 33530
rect 9330 33474 9382 33530
rect 7142 33250 9382 33474
rect 12446 33530 14686 33608
rect 12446 33474 12498 33530
rect 14322 33474 14686 33530
rect 12446 33250 14686 33474
rect 1480 33198 1838 33250
rect 1480 31062 1558 33198
rect 1614 31062 1838 33198
rect 1480 31010 1838 31062
tri 4471 31061 4611 31201 se
tri 4611 31131 4681 31201 sw
tri 4611 31061 4681 31131 nw
tri 6539 31131 6609 31201 se
tri 6609 31177 6633 31201 sw
tri 9891 31177 9915 31201 se
tri 6539 31061 6609 31131 ne
rect 6609 31061 6633 31177
tri 4420 31010 4471 31061 se
rect 0 30988 1240 31010
rect 0 30620 592 30988
rect 648 30620 1240 30988
tri 4331 30921 4420 31010 se
rect 4420 30921 4471 31010
tri 4471 30921 4611 31061 nw
tri 6609 31037 6633 31061 ne
tri 6633 31037 6773 31177 sw
tri 9775 31061 9891 31177 se
rect 9891 31061 9915 31177
tri 9915 31131 9985 31201 sw
tri 9915 31061 9985 31131 nw
tri 11843 31131 11913 31201 se
tri 11913 31177 11937 31201 sw
tri 11843 31061 11913 31131 ne
rect 11913 31061 11937 31177
tri 9751 31037 9775 31061 se
tri 6633 30921 6749 31037 ne
rect 6749 30921 6773 31037
tri 4191 30781 4331 30921 se
tri 4331 30781 4471 30921 nw
tri 6749 30897 6773 30921 ne
tri 6773 30897 6913 31037 sw
tri 9635 30921 9751 31037 se
rect 9751 30921 9775 31037
tri 9775 30921 9915 31061 nw
tri 11913 31037 11937 31061 ne
tri 11937 31037 12077 31177 sw
tri 11937 30921 12053 31037 ne
rect 12053 30921 12077 31037
tri 9611 30897 9635 30921 se
tri 6773 30781 6889 30897 ne
rect 6889 30781 6913 30897
tri 4051 30641 4191 30781 se
tri 4191 30641 4331 30781 nw
tri 6889 30757 6913 30781 ne
tri 6913 30757 7053 30897 sw
tri 9495 30781 9611 30897 se
rect 9611 30781 9635 30897
tri 9635 30781 9775 30921 nw
tri 12053 30897 12077 30921 ne
tri 12077 30897 12217 31037 sw
rect 15860 31010 15948 34424
rect 15284 30988 16524 31010
tri 12077 30781 12193 30897 ne
rect 12193 30781 12217 30897
tri 9471 30757 9495 30781 se
tri 6913 30641 7029 30757 ne
rect 7029 30641 7053 30757
rect 0 30598 1240 30620
tri 4008 30598 4051 30641 se
rect 576 28358 664 30598
tri 3911 30501 4008 30598 se
rect 4008 30501 4051 30598
tri 4051 30501 4191 30641 nw
tri 7029 30617 7053 30641 ne
tri 7053 30617 7193 30757 sw
tri 9355 30641 9471 30757 se
rect 9471 30641 9495 30757
tri 9495 30641 9635 30781 nw
tri 12193 30757 12217 30781 ne
tri 12217 30757 12357 30897 sw
tri 12217 30641 12333 30757 ne
rect 12333 30641 12357 30757
tri 9331 30617 9355 30641 se
tri 7053 30501 7169 30617 ne
rect 7169 30501 7193 30617
tri 3887 30477 3911 30501 se
rect 3911 30477 3957 30501
tri 3887 30407 3957 30477 ne
tri 3957 30407 4051 30501 nw
tri 7169 30477 7193 30501 ne
tri 7193 30477 7333 30617 sw
tri 9215 30501 9331 30617 se
rect 9331 30501 9355 30617
tri 9355 30501 9495 30641 nw
tri 12333 30617 12357 30641 ne
tri 12357 30617 12497 30757 sw
rect 15284 30620 15876 30988
rect 15932 30620 16524 30988
tri 12357 30501 12473 30617 ne
rect 12473 30501 12497 30617
tri 7193 30407 7263 30477 ne
tri 7263 30407 7333 30477 nw
tri 9191 30477 9215 30501 se
rect 9215 30477 9261 30501
tri 9191 30407 9261 30477 ne
tri 9261 30407 9355 30501 nw
tri 12473 30477 12497 30501 ne
tri 12497 30477 12637 30617 sw
rect 15284 30598 16524 30620
tri 12497 30407 12567 30477 ne
tri 12567 30407 12637 30477 nw
rect 14686 30546 15044 30598
tri 4471 28409 4611 28549 se
tri 4611 28479 4681 28549 sw
tri 4611 28409 4681 28479 nw
tri 6539 28479 6609 28549 se
tri 6609 28525 6633 28549 sw
tri 9891 28525 9915 28549 se
tri 6539 28409 6609 28479 ne
rect 6609 28409 6633 28525
tri 4420 28358 4471 28409 se
rect 0 28336 1240 28358
rect 0 27968 592 28336
rect 648 27968 1240 28336
tri 4331 28269 4420 28358 se
rect 4420 28269 4471 28358
tri 4471 28269 4611 28409 nw
tri 6609 28385 6633 28409 ne
tri 6633 28385 6773 28525 sw
tri 9775 28409 9891 28525 se
rect 9891 28409 9915 28525
tri 9915 28479 9985 28549 sw
tri 9915 28409 9985 28479 nw
tri 11843 28479 11913 28549 se
tri 11913 28525 11937 28549 sw
tri 11843 28409 11913 28479 ne
rect 11913 28409 11937 28525
tri 9751 28385 9775 28409 se
tri 6633 28269 6749 28385 ne
rect 6749 28269 6773 28385
tri 4191 28129 4331 28269 se
tri 4331 28129 4471 28269 nw
tri 6749 28245 6773 28269 ne
tri 6773 28245 6913 28385 sw
tri 9635 28269 9751 28385 se
rect 9751 28269 9775 28385
tri 9775 28269 9915 28409 nw
tri 11913 28385 11937 28409 ne
tri 11937 28385 12077 28525 sw
rect 14686 28410 14910 30546
rect 14966 28410 15044 30546
tri 11937 28269 12053 28385 ne
rect 12053 28269 12077 28385
tri 9611 28245 9635 28269 se
tri 6773 28129 6889 28245 ne
rect 6889 28129 6913 28245
tri 4051 27989 4191 28129 se
tri 4191 27989 4331 28129 nw
tri 6889 28105 6913 28129 ne
tri 6913 28105 7053 28245 sw
tri 9495 28129 9611 28245 se
rect 9611 28129 9635 28245
tri 9635 28129 9775 28269 nw
tri 12053 28245 12077 28269 ne
tri 12077 28245 12217 28385 sw
rect 14686 28358 15044 28410
rect 15860 28358 15948 30598
rect 15284 28336 16524 28358
tri 12077 28129 12193 28245 ne
rect 12193 28129 12217 28245
tri 9471 28105 9495 28129 se
tri 6913 27989 7029 28105 ne
rect 7029 27989 7053 28105
rect 0 27946 1240 27968
tri 4008 27946 4051 27989 se
rect 576 25706 664 27946
rect 1480 27894 1838 27946
rect 1480 25758 1558 27894
rect 1614 25758 1838 27894
tri 3911 27849 4008 27946 se
rect 4008 27849 4051 27946
tri 4051 27849 4191 27989 nw
tri 7029 27965 7053 27989 ne
tri 7053 27965 7193 28105 sw
tri 9355 27989 9471 28105 se
rect 9471 27989 9495 28105
tri 9495 27989 9635 28129 nw
tri 12193 28105 12217 28129 ne
tri 12217 28105 12357 28245 sw
tri 12217 27989 12333 28105 ne
rect 12333 27989 12357 28105
tri 9331 27965 9355 27989 se
tri 7053 27849 7169 27965 ne
rect 7169 27849 7193 27965
tri 3887 27825 3911 27849 se
rect 3911 27825 3957 27849
tri 3887 27755 3957 27825 ne
tri 3957 27755 4051 27849 nw
tri 7169 27825 7193 27849 ne
tri 7193 27825 7333 27965 sw
tri 9215 27849 9331 27965 se
rect 9331 27849 9355 27965
tri 9355 27849 9495 27989 nw
tri 12333 27965 12357 27989 ne
tri 12357 27965 12497 28105 sw
rect 15284 27968 15876 28336
rect 15932 27968 16524 28336
tri 12357 27849 12473 27965 ne
rect 12473 27849 12497 27965
tri 7193 27755 7263 27825 ne
tri 7263 27755 7333 27825 nw
tri 9191 27825 9215 27849 se
rect 9215 27825 9261 27849
tri 9191 27755 9261 27825 ne
tri 9261 27755 9355 27849 nw
tri 12473 27825 12497 27849 ne
tri 12497 27825 12637 27965 sw
rect 15284 27946 16524 27968
tri 12497 27755 12567 27825 ne
tri 12567 27755 12637 27825 nw
rect 1480 25706 1838 25758
tri 4471 25757 4611 25897 se
tri 4611 25827 4681 25897 sw
tri 4611 25757 4681 25827 nw
tri 6539 25827 6609 25897 se
tri 6609 25873 6633 25897 sw
tri 9891 25873 9915 25897 se
tri 6539 25757 6609 25827 ne
rect 6609 25757 6633 25873
tri 4420 25706 4471 25757 se
rect 0 25684 1240 25706
rect 0 25316 592 25684
rect 648 25316 1240 25684
tri 4331 25617 4420 25706 se
rect 4420 25617 4471 25706
tri 4471 25617 4611 25757 nw
tri 6609 25733 6633 25757 ne
tri 6633 25733 6773 25873 sw
tri 9775 25757 9891 25873 se
rect 9891 25757 9915 25873
tri 9915 25827 9985 25897 sw
tri 9915 25757 9985 25827 nw
tri 11843 25827 11913 25897 se
tri 11913 25873 11937 25897 sw
tri 11843 25757 11913 25827 ne
rect 11913 25757 11937 25873
tri 9751 25733 9775 25757 se
tri 6633 25617 6749 25733 ne
rect 6749 25617 6773 25733
tri 4191 25477 4331 25617 se
tri 4331 25477 4471 25617 nw
tri 6749 25593 6773 25617 ne
tri 6773 25593 6913 25733 sw
tri 9635 25617 9751 25733 se
rect 9751 25617 9775 25733
tri 9775 25617 9915 25757 nw
tri 11913 25733 11937 25757 ne
tri 11937 25733 12077 25873 sw
tri 11937 25617 12053 25733 ne
rect 12053 25617 12077 25733
tri 9611 25593 9635 25617 se
tri 6773 25477 6889 25593 ne
rect 6889 25477 6913 25593
tri 4051 25337 4191 25477 se
tri 4191 25337 4331 25477 nw
tri 6889 25453 6913 25477 ne
tri 6913 25453 7053 25593 sw
tri 9495 25477 9611 25593 se
rect 9611 25477 9635 25593
tri 9635 25477 9775 25617 nw
tri 12053 25593 12077 25617 ne
tri 12077 25593 12217 25733 sw
rect 15860 25706 15948 27946
rect 15284 25684 16524 25706
tri 12077 25477 12193 25593 ne
rect 12193 25477 12217 25593
tri 9471 25453 9495 25477 se
tri 6913 25337 7029 25453 ne
rect 7029 25337 7053 25453
rect 0 25294 1240 25316
tri 4008 25294 4051 25337 se
rect 576 23054 664 25294
tri 3911 25197 4008 25294 se
rect 4008 25197 4051 25294
tri 4051 25197 4191 25337 nw
tri 7029 25313 7053 25337 ne
tri 7053 25313 7193 25453 sw
tri 9355 25337 9471 25453 se
rect 9471 25337 9495 25453
tri 9495 25337 9635 25477 nw
tri 12193 25453 12217 25477 ne
tri 12217 25453 12357 25593 sw
tri 12217 25337 12333 25453 ne
rect 12333 25337 12357 25453
tri 9331 25313 9355 25337 se
tri 7053 25197 7169 25313 ne
rect 7169 25197 7193 25313
tri 3887 25173 3911 25197 se
rect 3911 25173 3957 25197
tri 3887 25103 3957 25173 ne
tri 3957 25103 4051 25197 nw
tri 7169 25173 7193 25197 ne
tri 7193 25173 7333 25313 sw
tri 9215 25197 9331 25313 se
rect 9331 25197 9355 25313
tri 9355 25197 9495 25337 nw
tri 12333 25313 12357 25337 ne
tri 12357 25313 12497 25453 sw
rect 15284 25316 15876 25684
rect 15932 25316 16524 25684
tri 12357 25197 12473 25313 ne
rect 12473 25197 12497 25313
tri 7193 25103 7263 25173 ne
tri 7263 25103 7333 25173 nw
tri 9191 25173 9215 25197 se
rect 9215 25173 9261 25197
tri 9191 25103 9261 25173 ne
tri 9261 25103 9355 25197 nw
tri 12473 25173 12497 25197 ne
tri 12497 25173 12637 25313 sw
rect 15284 25294 16524 25316
tri 12497 25103 12567 25173 ne
tri 12567 25103 12637 25173 nw
rect 14686 25242 15044 25294
rect 14686 23418 14910 25242
rect 14966 23418 15044 25242
tri 4471 23105 4611 23245 se
tri 4611 23175 4681 23245 sw
tri 4611 23105 4681 23175 nw
tri 6539 23175 6609 23245 se
tri 6609 23221 6633 23245 sw
tri 9891 23221 9915 23245 se
tri 6539 23105 6609 23175 ne
rect 6609 23105 6633 23221
tri 4420 23054 4471 23105 se
rect 0 23032 1240 23054
rect 0 22664 592 23032
rect 648 22664 1240 23032
tri 4331 22965 4420 23054 se
rect 4420 22965 4471 23054
tri 4471 22965 4611 23105 nw
tri 6609 23081 6633 23105 ne
tri 6633 23081 6773 23221 sw
tri 9775 23105 9891 23221 se
rect 9891 23105 9915 23221
tri 9915 23175 9985 23245 sw
tri 9915 23105 9985 23175 nw
tri 11843 23175 11913 23245 se
tri 11913 23221 11937 23245 sw
tri 11843 23105 11913 23175 ne
rect 11913 23105 11937 23221
tri 9751 23081 9775 23105 se
tri 6633 22965 6749 23081 ne
rect 6749 22965 6773 23081
tri 4191 22825 4331 22965 se
tri 4331 22825 4471 22965 nw
tri 6749 22941 6773 22965 ne
tri 6773 22941 6913 23081 sw
tri 9635 22965 9751 23081 se
rect 9751 22965 9775 23081
tri 9775 22965 9915 23105 nw
tri 11913 23081 11937 23105 ne
tri 11937 23081 12077 23221 sw
tri 11937 22965 12053 23081 ne
rect 12053 22965 12077 23081
tri 9611 22941 9635 22965 se
tri 6773 22825 6889 22941 ne
rect 6889 22825 6913 22941
tri 4051 22685 4191 22825 se
tri 4191 22685 4331 22825 nw
tri 6889 22801 6913 22825 ne
tri 6913 22801 7053 22941 sw
tri 9495 22825 9611 22941 se
rect 9611 22825 9635 22941
tri 9635 22825 9775 22965 nw
tri 12053 22941 12077 22965 ne
tri 12077 22941 12217 23081 sw
rect 14686 23054 15044 23418
rect 15860 23054 15948 25294
rect 15284 23032 16524 23054
tri 12077 22825 12193 22941 ne
rect 12193 22825 12217 22941
tri 9471 22801 9495 22825 se
tri 6913 22685 7029 22801 ne
rect 7029 22685 7053 22801
rect 0 22642 1240 22664
tri 4016 22650 4051 22685 se
rect 576 20402 664 22642
rect 1507 22590 1865 22650
rect 1507 20454 1558 22590
rect 1614 20454 1865 22590
tri 3911 22545 4016 22650 se
rect 4016 22545 4051 22650
tri 4051 22545 4191 22685 nw
tri 7029 22661 7053 22685 ne
tri 7053 22661 7193 22801 sw
tri 9355 22685 9471 22801 se
rect 9471 22685 9495 22801
tri 9495 22685 9635 22825 nw
tri 12193 22801 12217 22825 ne
tri 12217 22801 12357 22941 sw
tri 12217 22685 12333 22801 ne
rect 12333 22685 12357 22801
tri 9331 22661 9355 22685 se
tri 7053 22545 7169 22661 ne
rect 7169 22545 7193 22661
tri 3887 22521 3911 22545 se
rect 3911 22521 3957 22545
tri 3887 22451 3957 22521 ne
tri 3957 22451 4051 22545 nw
tri 7169 22521 7193 22545 ne
tri 7193 22521 7333 22661 sw
tri 9215 22545 9331 22661 se
rect 9331 22545 9355 22661
tri 9355 22545 9495 22685 nw
tri 12333 22661 12357 22685 ne
tri 12357 22661 12497 22801 sw
rect 15284 22664 15876 23032
rect 15932 22664 16524 23032
tri 12357 22545 12473 22661 ne
rect 12473 22545 12497 22661
tri 7193 22451 7263 22521 ne
tri 7263 22451 7333 22521 nw
tri 9191 22521 9215 22545 se
rect 9215 22521 9261 22545
tri 9191 22451 9261 22521 ne
tri 9261 22451 9355 22545 nw
tri 12473 22521 12497 22545 ne
tri 12497 22521 12637 22661 sw
rect 15284 22642 16524 22664
tri 12497 22451 12567 22521 ne
tri 12567 22451 12637 22521 nw
rect 1507 20410 1865 20454
tri 4471 20453 4611 20593 se
tri 4611 20523 4681 20593 sw
tri 4611 20453 4681 20523 nw
tri 6539 20523 6609 20593 se
tri 6609 20569 6633 20593 sw
tri 9891 20569 9915 20593 se
tri 6539 20453 6609 20523 ne
rect 6609 20453 6633 20569
tri 4428 20410 4471 20453 se
tri 4420 20402 4428 20410 se
rect 4428 20402 4471 20410
rect 0 20380 1240 20402
rect 0 20012 592 20380
rect 648 20012 1240 20380
tri 4331 20313 4420 20402 se
rect 4420 20313 4471 20402
tri 4471 20313 4611 20453 nw
tri 6609 20429 6633 20453 ne
tri 6633 20429 6773 20569 sw
tri 9775 20453 9891 20569 se
rect 9891 20453 9915 20569
tri 9915 20523 9985 20593 sw
tri 9915 20453 9985 20523 nw
tri 11843 20523 11913 20593 se
tri 11913 20569 11937 20593 sw
tri 11843 20453 11913 20523 ne
rect 11913 20453 11937 20569
tri 9751 20429 9775 20453 se
tri 6633 20313 6749 20429 ne
rect 6749 20313 6773 20429
tri 4191 20173 4331 20313 se
tri 4331 20173 4471 20313 nw
tri 6749 20289 6773 20313 ne
tri 6773 20289 6913 20429 sw
tri 9635 20313 9751 20429 se
rect 9751 20313 9775 20429
tri 9775 20313 9915 20453 nw
tri 11913 20429 11937 20453 ne
tri 11937 20429 12077 20569 sw
tri 11937 20313 12053 20429 ne
rect 12053 20313 12077 20429
tri 9611 20289 9635 20313 se
tri 6773 20173 6889 20289 ne
rect 6889 20173 6913 20289
tri 4051 20033 4191 20173 se
tri 4191 20033 4331 20173 nw
tri 6889 20149 6913 20173 ne
tri 6913 20149 7053 20289 sw
tri 9495 20173 9611 20289 se
rect 9611 20173 9635 20289
tri 9635 20173 9775 20313 nw
tri 12053 20289 12077 20313 ne
tri 12077 20289 12217 20429 sw
rect 15860 20402 15948 22642
rect 15284 20380 16524 20402
tri 12077 20173 12193 20289 ne
rect 12193 20173 12217 20289
tri 9471 20149 9495 20173 se
tri 6913 20033 7029 20149 ne
rect 7029 20033 7053 20149
rect 0 19990 1240 20012
tri 4008 19990 4051 20033 se
rect 576 17750 664 19990
tri 3911 19893 4008 19990 se
rect 4008 19893 4051 19990
tri 4051 19893 4191 20033 nw
tri 7029 20009 7053 20033 ne
tri 7053 20009 7193 20149 sw
tri 9355 20033 9471 20149 se
rect 9471 20033 9495 20149
tri 9495 20033 9635 20173 nw
tri 12193 20149 12217 20173 ne
tri 12217 20149 12357 20289 sw
tri 12217 20033 12333 20149 ne
rect 12333 20033 12357 20149
tri 9331 20009 9355 20033 se
tri 7053 19893 7169 20009 ne
rect 7169 19893 7193 20009
tri 3887 19869 3911 19893 se
rect 3911 19869 3957 19893
tri 3887 19799 3957 19869 ne
tri 3957 19799 4051 19893 nw
tri 7169 19869 7193 19893 ne
tri 7193 19869 7333 20009 sw
tri 9215 19893 9331 20009 se
rect 9331 19893 9355 20009
tri 9355 19893 9495 20033 nw
tri 12333 20009 12357 20033 ne
tri 12357 20009 12497 20149 sw
rect 15284 20012 15876 20380
rect 15932 20012 16524 20380
tri 12357 19893 12473 20009 ne
rect 12473 19893 12497 20009
tri 7193 19799 7263 19869 ne
tri 7263 19799 7333 19869 nw
tri 9191 19869 9215 19893 se
rect 9215 19869 9261 19893
tri 9191 19799 9261 19869 ne
tri 9261 19799 9355 19893 nw
tri 12473 19869 12497 19893 ne
tri 12497 19869 12637 20009 sw
rect 15284 19990 16524 20012
tri 12497 19799 12567 19869 ne
tri 12567 19799 12637 19869 nw
rect 14686 19938 15044 19990
tri 4471 17801 4611 17941 se
tri 4611 17871 4681 17941 sw
tri 4611 17801 4681 17871 nw
tri 6539 17871 6609 17941 se
tri 6609 17917 6633 17941 sw
tri 9891 17917 9915 17941 se
tri 6539 17801 6609 17871 ne
rect 6609 17801 6633 17917
tri 4420 17750 4471 17801 se
rect 0 17728 1240 17750
rect 0 17360 592 17728
rect 648 17360 1240 17728
tri 4331 17661 4420 17750 se
rect 4420 17661 4471 17750
tri 4471 17661 4611 17801 nw
tri 6609 17777 6633 17801 ne
tri 6633 17777 6773 17917 sw
tri 9775 17801 9891 17917 se
rect 9891 17801 9915 17917
tri 9915 17871 9985 17941 sw
tri 9915 17801 9985 17871 nw
tri 11843 17871 11913 17941 se
tri 11913 17917 11937 17941 sw
tri 11843 17801 11913 17871 ne
rect 11913 17801 11937 17917
tri 9751 17777 9775 17801 se
tri 6633 17661 6749 17777 ne
rect 6749 17661 6773 17777
tri 4191 17521 4331 17661 se
tri 4331 17521 4471 17661 nw
tri 6749 17637 6773 17661 ne
tri 6773 17637 6913 17777 sw
tri 9635 17661 9751 17777 se
rect 9751 17661 9775 17777
tri 9775 17661 9915 17801 nw
tri 11913 17777 11937 17801 ne
tri 11937 17777 12077 17917 sw
rect 14686 17802 14910 19938
rect 14966 17802 15044 19938
tri 11937 17661 12053 17777 ne
rect 12053 17661 12077 17777
tri 9611 17637 9635 17661 se
tri 6773 17521 6889 17637 ne
rect 6889 17521 6913 17637
tri 4051 17381 4191 17521 se
tri 4191 17381 4331 17521 nw
tri 6889 17497 6913 17521 ne
tri 6913 17497 7053 17637 sw
tri 9495 17521 9611 17637 se
rect 9611 17521 9635 17637
tri 9635 17521 9775 17661 nw
tri 12053 17637 12077 17661 ne
tri 12077 17637 12217 17777 sw
rect 14686 17750 15044 17802
rect 15860 17750 15948 19990
rect 15284 17728 16524 17750
tri 12077 17521 12193 17637 ne
rect 12193 17521 12217 17637
tri 9471 17497 9495 17521 se
tri 6913 17381 7029 17497 ne
rect 7029 17381 7053 17497
rect 0 17338 1240 17360
tri 4008 17338 4051 17381 se
rect 576 15098 664 17338
rect 1480 17286 1838 17338
rect 1480 15150 1558 17286
rect 1614 15150 1838 17286
tri 3911 17241 4008 17338 se
rect 4008 17241 4051 17338
tri 4051 17241 4191 17381 nw
tri 7029 17357 7053 17381 ne
tri 7053 17357 7193 17497 sw
tri 9355 17381 9471 17497 se
rect 9471 17381 9495 17497
tri 9495 17381 9635 17521 nw
tri 12193 17497 12217 17521 ne
tri 12217 17497 12357 17637 sw
tri 12217 17381 12333 17497 ne
rect 12333 17381 12357 17497
tri 9331 17357 9355 17381 se
tri 7053 17241 7169 17357 ne
rect 7169 17241 7193 17357
tri 3887 17217 3911 17241 se
rect 3911 17217 3957 17241
tri 3887 17147 3957 17217 ne
tri 3957 17147 4051 17241 nw
tri 7169 17217 7193 17241 ne
tri 7193 17217 7333 17357 sw
tri 9215 17241 9331 17357 se
rect 9331 17241 9355 17357
tri 9355 17241 9495 17381 nw
tri 12333 17357 12357 17381 ne
tri 12357 17357 12497 17497 sw
rect 15284 17360 15876 17728
rect 15932 17360 16524 17728
tri 12357 17241 12473 17357 ne
rect 12473 17241 12497 17357
tri 7193 17147 7263 17217 ne
tri 7263 17147 7333 17217 nw
tri 9191 17217 9215 17241 se
rect 9215 17217 9261 17241
tri 9191 17147 9261 17217 ne
tri 9261 17147 9355 17241 nw
tri 12473 17217 12497 17241 ne
tri 12497 17217 12637 17357 sw
rect 15284 17338 16524 17360
tri 12497 17147 12567 17217 ne
tri 12567 17147 12637 17217 nw
rect 1480 15098 1838 15150
tri 4471 15149 4611 15289 se
tri 4611 15219 4681 15289 sw
tri 4611 15149 4681 15219 nw
tri 6539 15219 6609 15289 se
tri 6609 15265 6633 15289 sw
tri 9891 15265 9915 15289 se
tri 6539 15149 6609 15219 ne
rect 6609 15149 6633 15265
tri 4420 15098 4471 15149 se
rect 0 15076 1240 15098
rect 0 14708 592 15076
rect 648 14708 1240 15076
tri 4331 15009 4420 15098 se
rect 4420 15009 4471 15098
tri 4471 15009 4611 15149 nw
tri 6609 15125 6633 15149 ne
tri 6633 15125 6773 15265 sw
tri 9775 15149 9891 15265 se
rect 9891 15149 9915 15265
tri 9915 15219 9985 15289 sw
tri 9915 15149 9985 15219 nw
tri 11843 15219 11913 15289 se
tri 11913 15265 11937 15289 sw
tri 11843 15149 11913 15219 ne
rect 11913 15149 11937 15265
tri 9751 15125 9775 15149 se
tri 6633 15009 6749 15125 ne
rect 6749 15009 6773 15125
tri 4191 14869 4331 15009 se
tri 4331 14869 4471 15009 nw
tri 6749 14985 6773 15009 ne
tri 6773 14985 6913 15125 sw
tri 9635 15009 9751 15125 se
rect 9751 15009 9775 15125
tri 9775 15009 9915 15149 nw
tri 11913 15125 11937 15149 ne
tri 11937 15125 12077 15265 sw
tri 11937 15009 12053 15125 ne
rect 12053 15009 12077 15125
tri 9611 14985 9635 15009 se
tri 6773 14869 6889 14985 ne
rect 6889 14869 6913 14985
tri 4051 14729 4191 14869 se
tri 4191 14729 4331 14869 nw
tri 6889 14845 6913 14869 ne
tri 6913 14845 7053 14985 sw
tri 9495 14869 9611 14985 se
rect 9611 14869 9635 14985
tri 9635 14869 9775 15009 nw
tri 12053 14985 12077 15009 ne
tri 12077 14985 12217 15125 sw
rect 15860 15098 15948 17338
rect 15284 15076 16524 15098
tri 12077 14869 12193 14985 ne
rect 12193 14869 12217 14985
tri 9471 14845 9495 14869 se
tri 6913 14729 7029 14845 ne
rect 7029 14729 7053 14845
rect 0 14686 1240 14708
tri 4008 14686 4051 14729 se
rect 576 12446 664 14686
tri 3911 14589 4008 14686 se
rect 4008 14589 4051 14686
tri 4051 14589 4191 14729 nw
tri 7029 14705 7053 14729 ne
tri 7053 14705 7193 14845 sw
tri 9355 14729 9471 14845 se
rect 9471 14729 9495 14845
tri 9495 14729 9635 14869 nw
tri 12193 14845 12217 14869 ne
tri 12217 14845 12357 14985 sw
tri 12217 14729 12333 14845 ne
rect 12333 14729 12357 14845
tri 9331 14705 9355 14729 se
tri 7053 14589 7169 14705 ne
rect 7169 14589 7193 14705
tri 3887 14565 3911 14589 se
rect 3911 14565 3957 14589
tri 3887 14495 3957 14565 ne
tri 3957 14495 4051 14589 nw
tri 7169 14565 7193 14589 ne
tri 7193 14565 7333 14705 sw
tri 9215 14589 9331 14705 se
rect 9331 14589 9355 14705
tri 9355 14589 9495 14729 nw
tri 12333 14705 12357 14729 ne
tri 12357 14705 12497 14845 sw
rect 15284 14708 15876 15076
rect 15932 14708 16524 15076
tri 12357 14589 12473 14705 ne
rect 12473 14589 12497 14705
tri 7193 14495 7263 14565 ne
tri 7263 14495 7333 14565 nw
tri 9191 14565 9215 14589 se
rect 9215 14565 9261 14589
tri 9191 14495 9261 14565 ne
tri 9261 14495 9355 14589 nw
tri 12473 14565 12497 14589 ne
tri 12497 14565 12637 14705 sw
rect 15284 14686 16524 14708
tri 12497 14495 12567 14565 ne
tri 12567 14495 12637 14565 nw
rect 14686 14634 15044 14686
rect 14686 12810 14910 14634
rect 14966 12810 15044 14634
tri 4471 12497 4611 12637 se
tri 4611 12567 4681 12637 sw
tri 4611 12497 4681 12567 nw
tri 6539 12567 6609 12637 se
tri 6609 12613 6633 12637 sw
tri 9891 12613 9915 12637 se
tri 6539 12497 6609 12567 ne
rect 6609 12497 6633 12613
tri 4420 12446 4471 12497 se
rect 0 12424 1240 12446
rect 0 12056 592 12424
rect 648 12056 1240 12424
tri 4331 12357 4420 12446 se
rect 4420 12357 4471 12446
tri 4471 12357 4611 12497 nw
tri 6609 12473 6633 12497 ne
tri 6633 12473 6773 12613 sw
tri 9775 12497 9891 12613 se
rect 9891 12497 9915 12613
tri 9915 12567 9985 12637 sw
tri 9915 12497 9985 12567 nw
tri 11843 12567 11913 12637 se
tri 11913 12613 11937 12637 sw
tri 11843 12497 11913 12567 ne
rect 11913 12497 11937 12613
tri 9751 12473 9775 12497 se
tri 6633 12357 6749 12473 ne
rect 6749 12357 6773 12473
tri 4191 12217 4331 12357 se
tri 4331 12217 4471 12357 nw
tri 6749 12333 6773 12357 ne
tri 6773 12333 6913 12473 sw
tri 9635 12357 9751 12473 se
rect 9751 12357 9775 12473
tri 9775 12357 9915 12497 nw
tri 11913 12473 11937 12497 ne
tri 11937 12473 12077 12613 sw
tri 11937 12357 12053 12473 ne
rect 12053 12357 12077 12473
tri 9611 12333 9635 12357 se
tri 6773 12217 6889 12333 ne
rect 6889 12217 6913 12333
tri 4051 12077 4191 12217 se
tri 4191 12077 4331 12217 nw
tri 6889 12193 6913 12217 ne
tri 6913 12193 7053 12333 sw
tri 9495 12217 9611 12333 se
rect 9611 12217 9635 12333
tri 9635 12217 9775 12357 nw
tri 12053 12333 12077 12357 ne
tri 12077 12333 12217 12473 sw
rect 14686 12446 15044 12810
rect 15860 12446 15948 14686
rect 15284 12424 16524 12446
tri 12077 12217 12193 12333 ne
rect 12193 12217 12217 12333
tri 9471 12193 9495 12217 se
tri 6913 12077 7029 12193 ne
rect 7029 12077 7053 12193
rect 0 12034 1240 12056
tri 4008 12034 4051 12077 se
rect 576 9794 664 12034
rect 1507 11982 1865 12034
rect 1507 9846 1558 11982
rect 1614 9846 1865 11982
tri 3911 11937 4008 12034 se
rect 4008 11937 4051 12034
tri 4051 11937 4191 12077 nw
tri 7029 12053 7053 12077 ne
tri 7053 12053 7193 12193 sw
tri 9355 12077 9471 12193 se
rect 9471 12077 9495 12193
tri 9495 12077 9635 12217 nw
tri 12193 12193 12217 12217 ne
tri 12217 12193 12357 12333 sw
tri 12217 12077 12333 12193 ne
rect 12333 12077 12357 12193
tri 9331 12053 9355 12077 se
tri 7053 11937 7169 12053 ne
rect 7169 11937 7193 12053
tri 3887 11913 3911 11937 se
rect 3911 11913 3957 11937
tri 3887 11843 3957 11913 ne
tri 3957 11843 4051 11937 nw
tri 7169 11913 7193 11937 ne
tri 7193 11913 7333 12053 sw
tri 9215 11937 9331 12053 se
rect 9331 11937 9355 12053
tri 9355 11937 9495 12077 nw
tri 12333 12053 12357 12077 ne
tri 12357 12053 12497 12193 sw
rect 15284 12056 15876 12424
rect 15932 12056 16524 12424
tri 12357 11937 12473 12053 ne
rect 12473 11937 12497 12053
tri 7193 11843 7263 11913 ne
tri 7263 11843 7333 11913 nw
tri 9191 11913 9215 11937 se
rect 9215 11913 9261 11937
tri 9191 11843 9261 11913 ne
tri 9261 11843 9355 11937 nw
tri 12473 11913 12497 11937 ne
tri 12497 11913 12637 12053 sw
rect 15284 12034 16524 12056
tri 12497 11843 12567 11913 ne
tri 12567 11843 12637 11913 nw
rect 1507 9794 1865 9846
tri 4471 9845 4611 9985 se
tri 4611 9915 4681 9985 sw
tri 4611 9845 4681 9915 nw
tri 6539 9915 6609 9985 se
tri 6609 9961 6633 9985 sw
tri 9891 9961 9915 9985 se
tri 6539 9845 6609 9915 ne
rect 6609 9845 6633 9961
tri 4420 9794 4471 9845 se
rect 0 9772 1240 9794
rect 0 9404 592 9772
rect 648 9404 1240 9772
tri 4331 9705 4420 9794 se
rect 4420 9705 4471 9794
tri 4471 9705 4611 9845 nw
tri 6609 9821 6633 9845 ne
tri 6633 9821 6773 9961 sw
tri 9775 9845 9891 9961 se
rect 9891 9845 9915 9961
tri 9915 9915 9985 9985 sw
tri 9915 9845 9985 9915 nw
tri 11843 9915 11913 9985 se
tri 11913 9961 11937 9985 sw
tri 11843 9845 11913 9915 ne
rect 11913 9845 11937 9961
tri 9751 9821 9775 9845 se
tri 6633 9705 6749 9821 ne
rect 6749 9705 6773 9821
tri 4191 9565 4331 9705 se
tri 4331 9565 4471 9705 nw
tri 6749 9681 6773 9705 ne
tri 6773 9681 6913 9821 sw
tri 9635 9705 9751 9821 se
rect 9751 9705 9775 9821
tri 9775 9705 9915 9845 nw
tri 11913 9821 11937 9845 ne
tri 11937 9821 12077 9961 sw
tri 11937 9705 12053 9821 ne
rect 12053 9705 12077 9821
tri 9611 9681 9635 9705 se
tri 6773 9565 6889 9681 ne
rect 6889 9565 6913 9681
tri 4051 9425 4191 9565 se
tri 4191 9425 4331 9565 nw
tri 6889 9541 6913 9565 ne
tri 6913 9541 7053 9681 sw
tri 9495 9565 9611 9681 se
rect 9611 9565 9635 9681
tri 9635 9565 9775 9705 nw
tri 12053 9681 12077 9705 ne
tri 12077 9681 12217 9821 sw
rect 15860 9794 15948 12034
rect 15284 9772 16524 9794
tri 12077 9565 12193 9681 ne
rect 12193 9565 12217 9681
tri 9471 9541 9495 9565 se
tri 6913 9425 7029 9541 ne
rect 7029 9425 7053 9541
rect 0 9382 1240 9404
tri 4008 9382 4051 9425 se
rect 576 7142 664 9382
tri 3911 9285 4008 9382 se
rect 4008 9285 4051 9382
tri 4051 9285 4191 9425 nw
tri 7029 9401 7053 9425 ne
tri 7053 9401 7193 9541 sw
tri 9355 9425 9471 9541 se
rect 9471 9425 9495 9541
tri 9495 9425 9635 9565 nw
tri 12193 9541 12217 9565 ne
tri 12217 9541 12357 9681 sw
tri 12217 9425 12333 9541 ne
rect 12333 9425 12357 9541
tri 9331 9401 9355 9425 se
tri 7053 9285 7169 9401 ne
rect 7169 9285 7193 9401
tri 3887 9261 3911 9285 se
rect 3911 9261 3957 9285
tri 3887 9191 3957 9261 ne
tri 3957 9191 4051 9285 nw
tri 7169 9261 7193 9285 ne
tri 7193 9261 7333 9401 sw
tri 9215 9285 9331 9401 se
rect 9331 9285 9355 9401
tri 9355 9285 9495 9425 nw
tri 12333 9401 12357 9425 ne
tri 12357 9401 12497 9541 sw
rect 15284 9404 15876 9772
rect 15932 9404 16524 9772
tri 12357 9285 12473 9401 ne
rect 12473 9285 12497 9401
tri 7193 9191 7263 9261 ne
tri 7263 9191 7333 9261 nw
tri 9191 9261 9215 9285 se
rect 9215 9261 9261 9285
tri 9191 9191 9261 9261 ne
tri 9261 9191 9355 9285 nw
tri 12473 9261 12497 9285 ne
tri 12497 9261 12637 9401 sw
rect 15284 9382 16524 9404
tri 12497 9191 12567 9261 ne
tri 12567 9191 12637 9261 nw
rect 14686 9330 15044 9382
tri 4471 7193 4611 7333 se
tri 4611 7263 4681 7333 sw
tri 4611 7193 4681 7263 nw
tri 6539 7263 6609 7333 se
tri 6609 7309 6633 7333 sw
tri 9891 7309 9915 7333 se
tri 6539 7193 6609 7263 ne
rect 6609 7193 6633 7309
tri 4420 7142 4471 7193 se
rect 0 7120 1240 7142
rect 0 6752 592 7120
rect 648 6752 1240 7120
tri 4331 7053 4420 7142 se
rect 4420 7053 4471 7142
tri 4471 7053 4611 7193 nw
tri 6609 7169 6633 7193 ne
tri 6633 7169 6773 7309 sw
tri 9775 7193 9891 7309 se
rect 9891 7193 9915 7309
tri 9915 7263 9985 7333 sw
tri 9915 7193 9985 7263 nw
tri 11843 7263 11913 7333 se
tri 11913 7309 11937 7333 sw
tri 11843 7193 11913 7263 ne
rect 11913 7193 11937 7309
tri 9751 7169 9775 7193 se
tri 6633 7053 6749 7169 ne
rect 6749 7053 6773 7169
tri 4191 6913 4331 7053 se
tri 4331 6913 4471 7053 nw
tri 6749 7029 6773 7053 ne
tri 6773 7029 6913 7169 sw
tri 9635 7053 9751 7169 se
rect 9751 7053 9775 7169
tri 9775 7053 9915 7193 nw
tri 11913 7169 11937 7193 ne
tri 11937 7169 12077 7309 sw
rect 14686 7194 14910 9330
rect 14966 7194 15044 9330
tri 11937 7053 12053 7169 ne
rect 12053 7053 12077 7169
tri 9611 7029 9635 7053 se
tri 6773 6913 6889 7029 ne
rect 6889 6913 6913 7029
tri 4051 6773 4191 6913 se
tri 4191 6773 4331 6913 nw
tri 6889 6889 6913 6913 ne
tri 6913 6889 7053 7029 sw
tri 9495 6913 9611 7029 se
rect 9611 6913 9635 7029
tri 9635 6913 9775 7053 nw
tri 12053 7029 12077 7053 ne
tri 12077 7029 12217 7169 sw
rect 14686 7142 15044 7194
rect 15860 7142 15948 9382
rect 15284 7120 16524 7142
tri 12077 6913 12193 7029 ne
rect 12193 6913 12217 7029
tri 9471 6889 9495 6913 se
tri 6913 6773 7029 6889 ne
rect 7029 6773 7053 6889
rect 0 6730 1240 6752
tri 4008 6730 4051 6773 se
rect 576 4490 664 6730
rect 1480 6678 1838 6730
rect 1480 4542 1558 6678
rect 1614 4542 1838 6678
tri 3911 6633 4008 6730 se
rect 4008 6633 4051 6730
tri 4051 6633 4191 6773 nw
tri 7029 6749 7053 6773 ne
tri 7053 6749 7193 6889 sw
tri 9355 6773 9471 6889 se
rect 9471 6773 9495 6889
tri 9495 6773 9635 6913 nw
tri 12193 6889 12217 6913 ne
tri 12217 6889 12357 7029 sw
tri 12217 6773 12333 6889 ne
rect 12333 6773 12357 6889
tri 9331 6749 9355 6773 se
tri 7053 6633 7169 6749 ne
rect 7169 6633 7193 6749
tri 3887 6609 3911 6633 se
rect 3911 6609 3957 6633
tri 3887 6539 3957 6609 ne
tri 3957 6539 4051 6633 nw
tri 7169 6609 7193 6633 ne
tri 7193 6609 7333 6749 sw
tri 9215 6633 9331 6749 se
rect 9331 6633 9355 6749
tri 9355 6633 9495 6773 nw
tri 12333 6749 12357 6773 ne
tri 12357 6749 12497 6889 sw
rect 15284 6752 15876 7120
rect 15932 6752 16524 7120
tri 12357 6633 12473 6749 ne
rect 12473 6633 12497 6749
tri 7193 6539 7263 6609 ne
tri 7263 6539 7333 6609 nw
tri 9191 6609 9215 6633 se
rect 9215 6609 9261 6633
tri 9191 6539 9261 6609 ne
tri 9261 6539 9355 6633 nw
tri 12473 6609 12497 6633 ne
tri 12497 6609 12637 6749 sw
rect 15284 6730 16524 6752
tri 12497 6539 12567 6609 ne
tri 12567 6539 12637 6609 nw
rect 1480 4490 1838 4542
tri 4471 4541 4611 4681 se
tri 4611 4611 4681 4681 sw
tri 4611 4541 4681 4611 nw
tri 6539 4611 6609 4681 se
tri 6609 4657 6633 4681 sw
tri 9891 4657 9915 4681 se
tri 6539 4541 6609 4611 ne
rect 6609 4541 6633 4657
tri 4420 4490 4471 4541 se
rect 0 4468 1240 4490
rect 0 4100 592 4468
rect 648 4100 1240 4468
tri 4331 4401 4420 4490 se
rect 4420 4401 4471 4490
tri 4471 4401 4611 4541 nw
tri 6609 4517 6633 4541 ne
tri 6633 4517 6773 4657 sw
tri 9775 4541 9891 4657 se
rect 9891 4541 9915 4657
tri 9915 4611 9985 4681 sw
tri 9915 4541 9985 4611 nw
tri 11843 4611 11913 4681 se
tri 11913 4657 11937 4681 sw
tri 11843 4541 11913 4611 ne
rect 11913 4541 11937 4657
tri 9751 4517 9775 4541 se
tri 6633 4401 6749 4517 ne
rect 6749 4401 6773 4517
tri 4191 4261 4331 4401 se
tri 4331 4261 4471 4401 nw
tri 6749 4377 6773 4401 ne
tri 6773 4377 6913 4517 sw
tri 9635 4401 9751 4517 se
rect 9751 4401 9775 4517
tri 9775 4401 9915 4541 nw
tri 11913 4517 11937 4541 ne
tri 11937 4517 12077 4657 sw
tri 11937 4401 12053 4517 ne
rect 12053 4401 12077 4517
tri 9611 4377 9635 4401 se
tri 6773 4261 6889 4377 ne
rect 6889 4261 6913 4377
tri 4051 4121 4191 4261 se
tri 4191 4121 4331 4261 nw
tri 6889 4237 6913 4261 ne
tri 6913 4237 7053 4377 sw
tri 9495 4261 9611 4377 se
rect 9611 4261 9635 4377
tri 9635 4261 9775 4401 nw
tri 12053 4377 12077 4401 ne
tri 12077 4377 12217 4517 sw
rect 15860 4490 15948 6730
rect 15284 4468 16524 4490
tri 12077 4261 12193 4377 ne
rect 12193 4261 12217 4377
tri 9471 4237 9495 4261 se
tri 6913 4121 7029 4237 ne
rect 7029 4121 7053 4237
rect 0 4078 1240 4100
tri 4008 4078 4051 4121 se
rect 576 664 664 4078
tri 3911 3981 4008 4078 se
rect 4008 3981 4051 4078
tri 4051 3981 4191 4121 nw
tri 7029 4097 7053 4121 ne
tri 7053 4097 7193 4237 sw
tri 9355 4121 9471 4237 se
rect 9471 4121 9495 4237
tri 9495 4121 9635 4261 nw
tri 12193 4237 12217 4261 ne
tri 12217 4237 12357 4377 sw
tri 12217 4121 12333 4237 ne
rect 12333 4121 12357 4237
tri 9331 4097 9355 4121 se
tri 7053 3981 7169 4097 ne
rect 7169 3981 7193 4097
tri 3887 3957 3911 3981 se
rect 3911 3957 3957 3981
tri 3887 3887 3957 3957 ne
tri 3957 3887 4051 3981 nw
tri 7169 3957 7193 3981 ne
tri 7193 3957 7333 4097 sw
tri 9215 3981 9331 4097 se
rect 9331 3981 9355 4097
tri 9355 3981 9495 4121 nw
tri 12333 4097 12357 4121 ne
tri 12357 4097 12497 4237 sw
rect 15284 4100 15876 4468
rect 15932 4100 16524 4468
tri 12357 3981 12473 4097 ne
rect 12473 3981 12497 4097
tri 7193 3887 7263 3957 ne
tri 7263 3887 7333 3957 nw
tri 9191 3957 9215 3981 se
rect 9215 3957 9261 3981
tri 9191 3887 9261 3957 ne
tri 9261 3887 9355 3981 nw
tri 12473 3957 12497 3981 ne
tri 12497 3957 12637 4097 sw
rect 15284 4078 16524 4100
tri 12497 3887 12567 3957 ne
tri 12567 3887 12637 3957 nw
rect 14686 4026 15044 4078
rect 14686 2202 14910 4026
rect 14966 2202 15044 4026
rect 14686 1838 15044 2202
rect 4490 1614 6730 1838
rect 4490 1558 4542 1614
rect 6678 1558 6730 1614
rect 4490 1480 6730 1558
rect 9794 1614 12034 1838
rect 9794 1558 9846 1614
rect 11982 1558 12034 1614
rect 9794 1480 12034 1558
rect 4078 664 4490 1240
rect 6730 664 7142 1240
rect 9382 664 9794 1240
rect 12034 664 12446 1240
rect 15860 664 15948 4078
rect 576 648 15948 664
rect 576 592 4100 648
rect 4468 592 6752 648
rect 7120 592 9404 648
rect 9772 592 12056 648
rect 12424 592 15948 648
rect 576 576 15948 592
rect 4078 0 4490 576
rect 6730 0 7142 576
rect 9382 0 9794 576
rect 12034 0 12446 576
<< via4 >>
rect 4100 34440 4468 34496
rect 6752 34440 7120 34496
rect 9404 34440 9772 34496
rect 12056 34440 12424 34496
rect 2202 33474 4026 33530
rect 7194 33474 9330 33530
rect 12498 33474 14322 33530
rect 1558 31062 1614 33198
rect 592 30620 648 30988
rect 15876 30620 15932 30988
rect 592 27968 648 28336
rect 14910 28410 14966 30546
rect 1558 25758 1614 27894
rect 15876 27968 15932 28336
rect 592 25316 648 25684
rect 15876 25316 15932 25684
rect 14910 23418 14966 25242
rect 592 22664 648 23032
rect 1558 20454 1614 22590
rect 15876 22664 15932 23032
rect 592 20012 648 20380
rect 15876 20012 15932 20380
rect 592 17360 648 17728
rect 14910 17802 14966 19938
rect 1558 15150 1614 17286
rect 15876 17360 15932 17728
rect 592 14708 648 15076
rect 15876 14708 15932 15076
rect 14910 12810 14966 14634
rect 592 12056 648 12424
rect 1558 9846 1614 11982
rect 15876 12056 15932 12424
rect 592 9404 648 9772
rect 15876 9404 15932 9772
rect 592 6752 648 7120
rect 14910 7194 14966 9330
rect 1558 4542 1614 6678
rect 15876 6752 15932 7120
rect 592 4100 648 4468
rect 15876 4100 15932 4468
rect 14910 2202 14966 4026
rect 4542 1558 6678 1614
rect 9846 1558 11982 1614
rect 4100 592 4468 648
rect 6752 592 7120 648
rect 9404 592 9772 648
rect 12056 592 12424 648
<< metal5 >>
rect 576 30988 664 34512
rect 576 30620 592 30988
rect 648 30620 664 30988
rect 576 28336 664 30620
rect 576 27968 592 28336
rect 648 27968 664 28336
rect 576 25684 664 27968
rect 576 25316 592 25684
rect 648 25316 664 25684
rect 576 23032 664 25316
rect 576 22664 592 23032
rect 648 22664 664 23032
rect 576 20380 664 22664
rect 576 20012 592 20380
rect 648 20012 664 20380
rect 576 17728 664 20012
rect 576 17360 592 17728
rect 648 17360 664 17728
rect 576 15076 664 17360
rect 576 14708 592 15076
rect 648 14708 664 15076
rect 576 12424 664 14708
rect 576 12056 592 12424
rect 648 12056 664 12424
rect 576 9772 664 12056
rect 576 9404 592 9772
rect 648 9404 664 9772
rect 576 7120 664 9404
rect 576 6752 592 7120
rect 648 6752 664 7120
rect 576 4468 664 6752
rect 576 4100 592 4468
rect 648 4100 664 4468
rect 576 664 664 4100
rect 1542 33198 1630 36415
rect 1542 31062 1558 33198
rect 1614 31062 1630 33198
rect 1542 27894 1630 31062
rect 1542 25758 1558 27894
rect 1614 25758 1630 27894
rect 1542 22590 1630 25758
rect 1542 20454 1558 22590
rect 1614 20454 1630 22590
rect 1542 17286 1630 20454
rect 1542 15150 1558 17286
rect 1614 15150 1630 17286
rect 1542 11982 1630 15150
rect 1542 9846 1558 11982
rect 1614 9846 1630 11982
rect 1542 6678 1630 9846
rect 1542 4542 1558 6678
rect 1614 4542 1630 6678
rect 1750 33130 1838 36415
rect 3958 34496 12566 34512
rect 3958 34440 4100 34496
rect 4468 34440 6752 34496
rect 7120 34440 9404 34496
rect 9772 34440 12056 34496
rect 12424 34440 12566 34496
rect 3958 34424 12566 34440
rect 2178 33530 14345 33546
rect 2178 33474 2202 33530
rect 4026 33474 7194 33530
rect 9330 33474 12498 33530
rect 14322 33474 14345 33530
rect 2178 33458 14345 33474
rect 14686 33338 14774 36415
rect 4610 33250 14774 33338
rect 4610 33130 6610 33250
rect 9914 33130 11914 33250
rect 1750 31130 1958 33130
tri 3887 31131 3957 31201 se
tri 3957 31131 4027 31201 sw
tri 7193 31131 7263 31201 se
tri 7263 31131 7333 31201 sw
tri 3887 31130 3888 31131 ne
rect 3888 31130 4027 31131
rect 1750 27826 1838 31130
tri 3888 30991 4027 31130 ne
tri 4027 30991 4167 31131 sw
tri 7169 31107 7193 31131 se
rect 7193 31107 7309 31131
tri 7309 31107 7333 31131 nw
tri 9191 31131 9261 31201 se
tri 9261 31131 9331 31201 sw
tri 12497 31131 12567 31201 se
tri 12567 31131 12637 31201 sw
tri 9191 31107 9215 31131 ne
rect 9215 31107 9331 31131
tri 7053 30991 7169 31107 se
tri 4027 30851 4167 30991 ne
tri 4167 30851 4307 30991 sw
tri 7029 30967 7053 30991 se
rect 7053 30967 7169 30991
tri 7169 30967 7309 31107 nw
tri 9215 30991 9331 31107 ne
tri 9331 30991 9471 31131 sw
tri 12473 31107 12497 31131 se
rect 12497 31107 12613 31131
tri 12613 31107 12637 31131 nw
tri 12357 30991 12473 31107 se
tri 9331 30967 9355 30991 ne
rect 9355 30967 9471 30991
tri 6913 30851 7029 30967 se
tri 4167 30711 4307 30851 ne
tri 4307 30711 4447 30851 sw
tri 6889 30827 6913 30851 se
rect 6913 30827 7029 30851
tri 7029 30827 7169 30967 nw
tri 9355 30851 9471 30967 ne
tri 9471 30851 9611 30991 sw
tri 12333 30967 12357 30991 se
rect 12357 30967 12473 30991
tri 12473 30967 12613 31107 nw
tri 12217 30851 12333 30967 se
tri 9471 30827 9495 30851 ne
rect 9495 30827 9611 30851
tri 6773 30711 6889 30827 se
tri 4307 30571 4447 30711 ne
tri 4447 30571 4587 30711 sw
tri 6749 30687 6773 30711 se
rect 6773 30687 6889 30711
tri 6889 30687 7029 30827 nw
tri 9495 30711 9611 30827 ne
tri 9611 30711 9751 30851 sw
tri 12193 30827 12217 30851 se
rect 12217 30827 12333 30851
tri 12333 30827 12473 30967 nw
tri 12077 30711 12193 30827 se
tri 9611 30687 9635 30711 ne
rect 9635 30687 9751 30711
tri 6633 30571 6749 30687 se
tri 4447 30431 4587 30571 ne
tri 4587 30477 4681 30571 sw
tri 6609 30547 6633 30571 se
rect 6633 30547 6749 30571
tri 6749 30547 6889 30687 nw
tri 9635 30571 9751 30687 ne
tri 9751 30571 9891 30711 sw
tri 12053 30687 12077 30711 se
rect 12077 30687 12193 30711
tri 12193 30687 12333 30827 nw
tri 11937 30571 12053 30687 se
tri 9751 30547 9775 30571 ne
rect 9775 30547 9891 30571
rect 4587 30431 4611 30477
tri 4587 30407 4611 30431 ne
tri 4611 30407 4681 30477 nw
tri 6539 30477 6609 30547 se
tri 6539 30407 6609 30477 ne
tri 6609 30407 6749 30547 nw
tri 9775 30431 9891 30547 ne
tri 9891 30477 9985 30571 sw
tri 11913 30547 11937 30571 se
rect 11937 30547 12053 30571
tri 12053 30547 12193 30687 nw
rect 9891 30431 9915 30477
tri 9891 30407 9915 30431 ne
tri 9915 30407 9985 30477 nw
tri 11843 30477 11913 30547 se
tri 11843 30407 11913 30477 ne
tri 11913 30407 12053 30547 nw
rect 14686 30478 14774 33250
tri 3887 28479 3957 28549 se
tri 3957 28479 4027 28549 sw
tri 7193 28479 7263 28549 se
tri 7263 28479 7333 28549 sw
tri 3887 28339 4027 28479 ne
tri 4027 28339 4167 28479 sw
tri 7169 28455 7193 28479 se
rect 7193 28455 7309 28479
tri 7309 28455 7333 28479 nw
tri 9191 28479 9261 28549 se
tri 9261 28479 9331 28549 sw
tri 12497 28479 12567 28549 se
tri 12567 28479 12637 28549 sw
tri 9191 28455 9215 28479 ne
rect 9215 28455 9331 28479
tri 7053 28339 7169 28455 se
tri 4027 28199 4167 28339 ne
tri 4167 28199 4307 28339 sw
tri 7029 28315 7053 28339 se
rect 7053 28315 7169 28339
tri 7169 28315 7309 28455 nw
tri 9215 28339 9331 28455 ne
tri 9331 28339 9471 28479 sw
tri 12473 28455 12497 28479 se
rect 12497 28455 12613 28479
tri 12613 28455 12637 28479 nw
rect 14566 28478 14774 30478
tri 12357 28339 12473 28455 se
tri 9331 28315 9355 28339 ne
rect 9355 28315 9471 28339
tri 6913 28199 7029 28315 se
tri 4167 28059 4307 28199 ne
tri 4307 28059 4447 28199 sw
tri 6889 28175 6913 28199 se
rect 6913 28175 7029 28199
tri 7029 28175 7169 28315 nw
tri 9355 28199 9471 28315 ne
tri 9471 28199 9611 28339 sw
tri 12333 28315 12357 28339 se
rect 12357 28315 12473 28339
tri 12473 28315 12613 28455 nw
tri 12217 28199 12333 28315 se
tri 9471 28175 9495 28199 ne
rect 9495 28175 9611 28199
tri 6773 28059 6889 28175 se
tri 4307 27919 4447 28059 ne
tri 4447 27919 4587 28059 sw
tri 6749 28035 6773 28059 se
rect 6773 28035 6889 28059
tri 6889 28035 7029 28175 nw
tri 9495 28059 9611 28175 ne
tri 9611 28059 9751 28199 sw
tri 12193 28175 12217 28199 se
rect 12217 28175 12333 28199
tri 12333 28175 12473 28315 nw
tri 12077 28059 12193 28175 se
tri 9611 28035 9635 28059 ne
rect 9635 28035 9751 28059
tri 6633 27919 6749 28035 se
tri 4447 27826 4540 27919 ne
rect 4540 27826 4587 27919
rect 1750 25826 1958 27826
tri 4540 27779 4587 27826 ne
tri 4587 27825 4681 27919 sw
tri 6609 27895 6633 27919 se
rect 6633 27895 6749 27919
tri 6749 27895 6889 28035 nw
tri 9635 27919 9751 28035 ne
tri 9751 27919 9891 28059 sw
tri 12053 28035 12077 28059 se
rect 12077 28035 12193 28059
tri 12193 28035 12333 28175 nw
tri 11937 27919 12053 28035 se
tri 9751 27895 9775 27919 ne
rect 9775 27895 9891 27919
rect 4587 27779 4611 27825
tri 4587 27755 4611 27779 ne
tri 4611 27755 4681 27825 nw
tri 6539 27825 6609 27895 se
tri 6539 27755 6609 27825 ne
tri 6609 27755 6749 27895 nw
tri 9775 27779 9891 27895 ne
tri 9891 27825 9985 27919 sw
tri 11913 27895 11937 27919 se
rect 11937 27895 12053 27919
tri 12053 27895 12193 28035 nw
rect 9891 27779 9915 27825
tri 9891 27755 9915 27779 ne
tri 9915 27755 9985 27825 nw
tri 11843 27825 11913 27895 se
tri 11843 27755 11913 27825 ne
tri 11913 27755 12053 27895 nw
tri 3887 25827 3957 25897 se
tri 3957 25827 4027 25897 sw
tri 7193 25827 7263 25897 se
tri 7263 25827 7333 25897 sw
tri 3887 25826 3888 25827 ne
rect 3888 25826 4027 25827
rect 1750 22522 1838 25826
tri 3888 25687 4027 25826 ne
tri 4027 25687 4167 25827 sw
tri 7169 25803 7193 25827 se
rect 7193 25803 7309 25827
tri 7309 25803 7333 25827 nw
tri 9191 25827 9261 25897 se
tri 9261 25827 9331 25897 sw
tri 12497 25827 12567 25897 se
tri 12567 25827 12637 25897 sw
tri 9191 25803 9215 25827 ne
rect 9215 25803 9331 25827
tri 7053 25687 7169 25803 se
tri 4027 25547 4167 25687 ne
tri 4167 25547 4307 25687 sw
tri 7029 25663 7053 25687 se
rect 7053 25663 7169 25687
tri 7169 25663 7309 25803 nw
tri 9215 25687 9331 25803 ne
tri 9331 25687 9471 25827 sw
tri 12473 25803 12497 25827 se
rect 12497 25803 12613 25827
tri 12613 25803 12637 25827 nw
tri 12357 25687 12473 25803 se
tri 9331 25663 9355 25687 ne
rect 9355 25663 9471 25687
tri 6913 25547 7029 25663 se
tri 4167 25407 4307 25547 ne
tri 4307 25407 4447 25547 sw
tri 6889 25523 6913 25547 se
rect 6913 25523 7029 25547
tri 7029 25523 7169 25663 nw
tri 9355 25547 9471 25663 ne
tri 9471 25547 9611 25687 sw
tri 12333 25663 12357 25687 se
rect 12357 25663 12473 25687
tri 12473 25663 12613 25803 nw
tri 12217 25547 12333 25663 se
tri 9471 25523 9495 25547 ne
rect 9495 25523 9611 25547
tri 6773 25407 6889 25523 se
tri 4307 25267 4447 25407 ne
tri 4447 25267 4587 25407 sw
tri 6749 25383 6773 25407 se
rect 6773 25383 6889 25407
tri 6889 25383 7029 25523 nw
tri 9495 25407 9611 25523 ne
tri 9611 25407 9751 25547 sw
tri 12193 25523 12217 25547 se
rect 12217 25523 12333 25547
tri 12333 25523 12473 25663 nw
tri 12077 25407 12193 25523 se
tri 9611 25383 9635 25407 ne
rect 9635 25383 9751 25407
tri 6633 25267 6749 25383 se
tri 4447 25127 4587 25267 ne
tri 4587 25173 4681 25267 sw
tri 6609 25243 6633 25267 se
rect 6633 25243 6749 25267
tri 6749 25243 6889 25383 nw
tri 9635 25267 9751 25383 ne
tri 9751 25267 9891 25407 sw
tri 12053 25383 12077 25407 se
rect 12077 25383 12193 25407
tri 12193 25383 12333 25523 nw
tri 11937 25267 12053 25383 se
tri 9751 25243 9775 25267 ne
rect 9775 25243 9891 25267
rect 4587 25127 4611 25173
tri 4587 25103 4611 25127 ne
tri 4611 25103 4681 25173 nw
tri 6539 25173 6609 25243 se
tri 6539 25103 6609 25173 ne
tri 6609 25103 6749 25243 nw
tri 9775 25127 9891 25243 ne
tri 9891 25173 9985 25267 sw
tri 11913 25243 11937 25267 se
rect 11937 25243 12053 25267
tri 12053 25243 12193 25383 nw
rect 9891 25127 9915 25173
tri 9891 25103 9915 25127 ne
tri 9915 25103 9985 25173 nw
tri 11843 25173 11913 25243 se
tri 11843 25103 11913 25173 ne
tri 11913 25103 12053 25243 nw
rect 14686 25174 14774 28478
tri 3887 23175 3957 23245 se
tri 3957 23175 4027 23245 sw
tri 7193 23175 7263 23245 se
tri 7263 23175 7333 23245 sw
tri 3887 23035 4027 23175 ne
tri 4027 23035 4167 23175 sw
tri 7169 23151 7193 23175 se
rect 7193 23151 7309 23175
tri 7309 23151 7333 23175 nw
tri 9191 23175 9261 23245 se
tri 9261 23175 9331 23245 sw
tri 12497 23175 12567 23245 se
tri 12567 23175 12637 23245 sw
tri 9191 23151 9215 23175 ne
rect 9215 23151 9331 23175
tri 7053 23035 7169 23151 se
tri 4027 22895 4167 23035 ne
tri 4167 22895 4307 23035 sw
tri 7029 23011 7053 23035 se
rect 7053 23011 7169 23035
tri 7169 23011 7309 23151 nw
tri 9215 23035 9331 23151 ne
tri 9331 23035 9471 23175 sw
tri 12473 23151 12497 23175 se
rect 12497 23151 12613 23175
tri 12613 23151 12637 23175 nw
rect 14566 23174 14774 25174
tri 12357 23035 12473 23151 se
tri 9331 23011 9355 23035 ne
rect 9355 23011 9471 23035
tri 6913 22895 7029 23011 se
tri 4167 22755 4307 22895 ne
tri 4307 22755 4447 22895 sw
tri 6889 22871 6913 22895 se
rect 6913 22871 7029 22895
tri 7029 22871 7169 23011 nw
tri 9355 22895 9471 23011 ne
tri 9471 22895 9611 23035 sw
tri 12333 23011 12357 23035 se
rect 12357 23011 12473 23035
tri 12473 23011 12613 23151 nw
tri 12217 22895 12333 23011 se
tri 9471 22871 9495 22895 ne
rect 9495 22871 9611 22895
tri 6773 22755 6889 22871 se
tri 4307 22615 4447 22755 ne
tri 4447 22615 4587 22755 sw
tri 6749 22731 6773 22755 se
rect 6773 22731 6889 22755
tri 6889 22731 7029 22871 nw
tri 9495 22755 9611 22871 ne
tri 9611 22755 9751 22895 sw
tri 12193 22871 12217 22895 se
rect 12217 22871 12333 22895
tri 12333 22871 12473 23011 nw
tri 12077 22755 12193 22871 se
tri 9611 22731 9635 22755 ne
rect 9635 22731 9751 22755
tri 6633 22615 6749 22731 se
tri 4447 22522 4540 22615 ne
rect 4540 22522 4587 22615
rect 1750 20522 1958 22522
tri 4540 22475 4587 22522 ne
tri 4587 22521 4681 22615 sw
tri 6609 22591 6633 22615 se
rect 6633 22591 6749 22615
tri 6749 22591 6889 22731 nw
tri 9635 22615 9751 22731 ne
tri 9751 22615 9891 22755 sw
tri 12053 22731 12077 22755 se
rect 12077 22731 12193 22755
tri 12193 22731 12333 22871 nw
tri 11937 22615 12053 22731 se
tri 9751 22591 9775 22615 ne
rect 9775 22591 9891 22615
rect 4587 22475 4611 22521
tri 4587 22451 4611 22475 ne
tri 4611 22451 4681 22521 nw
tri 6539 22521 6609 22591 se
tri 6539 22451 6609 22521 ne
tri 6609 22451 6749 22591 nw
tri 9775 22475 9891 22591 ne
tri 9891 22521 9985 22615 sw
tri 11913 22591 11937 22615 se
rect 11937 22591 12053 22615
tri 12053 22591 12193 22731 nw
rect 9891 22475 9915 22521
tri 9891 22451 9915 22475 ne
tri 9915 22451 9985 22521 nw
tri 11843 22521 11913 22591 se
tri 11843 22451 11913 22521 ne
tri 11913 22451 12053 22591 nw
tri 3887 20523 3957 20593 se
tri 3957 20523 4027 20593 sw
tri 7193 20523 7263 20593 se
tri 7263 20523 7333 20593 sw
tri 3887 20522 3888 20523 ne
rect 3888 20522 4027 20523
rect 1750 17218 1838 20522
tri 3888 20383 4027 20522 ne
tri 4027 20383 4167 20523 sw
tri 7169 20499 7193 20523 se
rect 7193 20499 7309 20523
tri 7309 20499 7333 20523 nw
tri 9191 20523 9261 20593 se
tri 9261 20523 9331 20593 sw
tri 12497 20523 12567 20593 se
tri 12567 20523 12637 20593 sw
tri 9191 20499 9215 20523 ne
rect 9215 20499 9331 20523
tri 7053 20383 7169 20499 se
tri 4027 20243 4167 20383 ne
tri 4167 20243 4307 20383 sw
tri 7029 20359 7053 20383 se
rect 7053 20359 7169 20383
tri 7169 20359 7309 20499 nw
tri 9215 20383 9331 20499 ne
tri 9331 20383 9471 20523 sw
tri 12473 20499 12497 20523 se
rect 12497 20499 12613 20523
tri 12613 20499 12637 20523 nw
tri 12357 20383 12473 20499 se
tri 9331 20359 9355 20383 ne
rect 9355 20359 9471 20383
tri 6913 20243 7029 20359 se
tri 4167 20103 4307 20243 ne
tri 4307 20103 4447 20243 sw
tri 6889 20219 6913 20243 se
rect 6913 20219 7029 20243
tri 7029 20219 7169 20359 nw
tri 9355 20243 9471 20359 ne
tri 9471 20243 9611 20383 sw
tri 12333 20359 12357 20383 se
rect 12357 20359 12473 20383
tri 12473 20359 12613 20499 nw
tri 12217 20243 12333 20359 se
tri 9471 20219 9495 20243 ne
rect 9495 20219 9611 20243
tri 6773 20103 6889 20219 se
tri 4307 19963 4447 20103 ne
tri 4447 19963 4587 20103 sw
tri 6749 20079 6773 20103 se
rect 6773 20079 6889 20103
tri 6889 20079 7029 20219 nw
tri 9495 20103 9611 20219 ne
tri 9611 20103 9751 20243 sw
tri 12193 20219 12217 20243 se
rect 12217 20219 12333 20243
tri 12333 20219 12473 20359 nw
tri 12077 20103 12193 20219 se
tri 9611 20079 9635 20103 ne
rect 9635 20079 9751 20103
tri 6633 19963 6749 20079 se
tri 4447 19823 4587 19963 ne
tri 4587 19869 4681 19963 sw
tri 6609 19939 6633 19963 se
rect 6633 19939 6749 19963
tri 6749 19939 6889 20079 nw
tri 9635 19963 9751 20079 ne
tri 9751 19963 9891 20103 sw
tri 12053 20079 12077 20103 se
rect 12077 20079 12193 20103
tri 12193 20079 12333 20219 nw
tri 11937 19963 12053 20079 se
tri 9751 19939 9775 19963 ne
rect 9775 19939 9891 19963
rect 4587 19823 4611 19869
tri 4587 19799 4611 19823 ne
tri 4611 19799 4681 19869 nw
tri 6539 19869 6609 19939 se
tri 6539 19799 6609 19869 ne
tri 6609 19799 6749 19939 nw
tri 9775 19823 9891 19939 ne
tri 9891 19869 9985 19963 sw
tri 11913 19939 11937 19963 se
rect 11937 19939 12053 19963
tri 12053 19939 12193 20079 nw
rect 9891 19823 9915 19869
tri 9891 19799 9915 19823 ne
tri 9915 19799 9985 19869 nw
tri 11843 19869 11913 19939 se
tri 11843 19799 11913 19869 ne
tri 11913 19799 12053 19939 nw
rect 14686 19870 14774 23174
tri 3887 17871 3957 17941 se
tri 3957 17871 4027 17941 sw
tri 7193 17871 7263 17941 se
tri 7263 17871 7333 17941 sw
tri 3887 17731 4027 17871 ne
tri 4027 17731 4167 17871 sw
tri 7169 17847 7193 17871 se
rect 7193 17847 7309 17871
tri 7309 17847 7333 17871 nw
tri 9191 17871 9261 17941 se
tri 9261 17871 9331 17941 sw
tri 12497 17871 12567 17941 se
tri 12567 17871 12637 17941 sw
tri 9191 17847 9215 17871 ne
rect 9215 17847 9331 17871
tri 7053 17731 7169 17847 se
tri 4027 17591 4167 17731 ne
tri 4167 17591 4307 17731 sw
tri 7029 17707 7053 17731 se
rect 7053 17707 7169 17731
tri 7169 17707 7309 17847 nw
tri 9215 17731 9331 17847 ne
tri 9331 17731 9471 17871 sw
tri 12473 17847 12497 17871 se
rect 12497 17847 12613 17871
tri 12613 17847 12637 17871 nw
rect 14566 17870 14774 19870
tri 12357 17731 12473 17847 se
tri 9331 17707 9355 17731 ne
rect 9355 17707 9471 17731
tri 6913 17591 7029 17707 se
tri 4167 17451 4307 17591 ne
tri 4307 17451 4447 17591 sw
tri 6889 17567 6913 17591 se
rect 6913 17567 7029 17591
tri 7029 17567 7169 17707 nw
tri 9355 17591 9471 17707 ne
tri 9471 17591 9611 17731 sw
tri 12333 17707 12357 17731 se
rect 12357 17707 12473 17731
tri 12473 17707 12613 17847 nw
tri 12217 17591 12333 17707 se
tri 9471 17567 9495 17591 ne
rect 9495 17567 9611 17591
tri 6773 17451 6889 17567 se
tri 4307 17311 4447 17451 ne
tri 4447 17311 4587 17451 sw
tri 6749 17427 6773 17451 se
rect 6773 17427 6889 17451
tri 6889 17427 7029 17567 nw
tri 9495 17451 9611 17567 ne
tri 9611 17451 9751 17591 sw
tri 12193 17567 12217 17591 se
rect 12217 17567 12333 17591
tri 12333 17567 12473 17707 nw
tri 12077 17451 12193 17567 se
tri 9611 17427 9635 17451 ne
rect 9635 17427 9751 17451
tri 6633 17311 6749 17427 se
tri 4447 17218 4540 17311 ne
rect 4540 17218 4587 17311
rect 1750 15218 1958 17218
tri 4540 17171 4587 17218 ne
tri 4587 17217 4681 17311 sw
tri 6609 17287 6633 17311 se
rect 6633 17287 6749 17311
tri 6749 17287 6889 17427 nw
tri 9635 17311 9751 17427 ne
tri 9751 17311 9891 17451 sw
tri 12053 17427 12077 17451 se
rect 12077 17427 12193 17451
tri 12193 17427 12333 17567 nw
tri 11937 17311 12053 17427 se
tri 9751 17287 9775 17311 ne
rect 9775 17287 9891 17311
rect 4587 17171 4611 17217
tri 4587 17147 4611 17171 ne
tri 4611 17147 4681 17217 nw
tri 6539 17217 6609 17287 se
tri 6539 17147 6609 17217 ne
tri 6609 17147 6749 17287 nw
tri 9775 17171 9891 17287 ne
tri 9891 17217 9985 17311 sw
tri 11913 17287 11937 17311 se
rect 11937 17287 12053 17311
tri 12053 17287 12193 17427 nw
rect 9891 17171 9915 17217
tri 9891 17147 9915 17171 ne
tri 9915 17147 9985 17217 nw
tri 11843 17217 11913 17287 se
tri 11843 17147 11913 17217 ne
tri 11913 17147 12053 17287 nw
tri 3887 15219 3957 15289 se
tri 3957 15219 4027 15289 sw
tri 7193 15219 7263 15289 se
tri 7263 15219 7333 15289 sw
tri 3887 15218 3888 15219 ne
rect 3888 15218 4027 15219
rect 1750 11914 1838 15218
tri 3888 15079 4027 15218 ne
tri 4027 15079 4167 15219 sw
tri 7169 15195 7193 15219 se
rect 7193 15195 7309 15219
tri 7309 15195 7333 15219 nw
tri 9191 15219 9261 15289 se
tri 9261 15219 9331 15289 sw
tri 12497 15219 12567 15289 se
tri 12567 15219 12637 15289 sw
tri 9191 15195 9215 15219 ne
rect 9215 15195 9331 15219
tri 7053 15079 7169 15195 se
tri 4027 14939 4167 15079 ne
tri 4167 14939 4307 15079 sw
tri 7029 15055 7053 15079 se
rect 7053 15055 7169 15079
tri 7169 15055 7309 15195 nw
tri 9215 15079 9331 15195 ne
tri 9331 15079 9471 15219 sw
tri 12473 15195 12497 15219 se
rect 12497 15195 12613 15219
tri 12613 15195 12637 15219 nw
tri 12357 15079 12473 15195 se
tri 9331 15055 9355 15079 ne
rect 9355 15055 9471 15079
tri 6913 14939 7029 15055 se
tri 4167 14799 4307 14939 ne
tri 4307 14799 4447 14939 sw
tri 6889 14915 6913 14939 se
rect 6913 14915 7029 14939
tri 7029 14915 7169 15055 nw
tri 9355 14939 9471 15055 ne
tri 9471 14939 9611 15079 sw
tri 12333 15055 12357 15079 se
rect 12357 15055 12473 15079
tri 12473 15055 12613 15195 nw
tri 12217 14939 12333 15055 se
tri 9471 14915 9495 14939 ne
rect 9495 14915 9611 14939
tri 6773 14799 6889 14915 se
tri 4307 14659 4447 14799 ne
tri 4447 14659 4587 14799 sw
tri 6749 14775 6773 14799 se
rect 6773 14775 6889 14799
tri 6889 14775 7029 14915 nw
tri 9495 14799 9611 14915 ne
tri 9611 14799 9751 14939 sw
tri 12193 14915 12217 14939 se
rect 12217 14915 12333 14939
tri 12333 14915 12473 15055 nw
tri 12077 14799 12193 14915 se
tri 9611 14775 9635 14799 ne
rect 9635 14775 9751 14799
tri 6633 14659 6749 14775 se
tri 4447 14519 4587 14659 ne
tri 4587 14565 4681 14659 sw
tri 6609 14635 6633 14659 se
rect 6633 14635 6749 14659
tri 6749 14635 6889 14775 nw
tri 9635 14659 9751 14775 ne
tri 9751 14659 9891 14799 sw
tri 12053 14775 12077 14799 se
rect 12077 14775 12193 14799
tri 12193 14775 12333 14915 nw
tri 11937 14659 12053 14775 se
tri 9751 14635 9775 14659 ne
rect 9775 14635 9891 14659
rect 4587 14519 4611 14565
tri 4587 14495 4611 14519 ne
tri 4611 14495 4681 14565 nw
tri 6539 14565 6609 14635 se
tri 6539 14495 6609 14565 ne
tri 6609 14495 6749 14635 nw
tri 9775 14519 9891 14635 ne
tri 9891 14565 9985 14659 sw
tri 11913 14635 11937 14659 se
rect 11937 14635 12053 14659
tri 12053 14635 12193 14775 nw
rect 9891 14519 9915 14565
tri 9891 14495 9915 14519 ne
tri 9915 14495 9985 14565 nw
tri 11843 14565 11913 14635 se
tri 11843 14495 11913 14565 ne
tri 11913 14495 12053 14635 nw
rect 14686 14566 14774 17870
tri 3887 12567 3957 12637 se
tri 3957 12567 4027 12637 sw
tri 7193 12567 7263 12637 se
tri 7263 12567 7333 12637 sw
tri 3887 12427 4027 12567 ne
tri 4027 12427 4167 12567 sw
tri 7169 12543 7193 12567 se
rect 7193 12543 7309 12567
tri 7309 12543 7333 12567 nw
tri 9191 12567 9261 12637 se
tri 9261 12567 9331 12637 sw
tri 12497 12567 12567 12637 se
tri 12567 12567 12637 12637 sw
tri 9191 12543 9215 12567 ne
rect 9215 12543 9331 12567
tri 7053 12427 7169 12543 se
tri 4027 12287 4167 12427 ne
tri 4167 12287 4307 12427 sw
tri 7029 12403 7053 12427 se
rect 7053 12403 7169 12427
tri 7169 12403 7309 12543 nw
tri 9215 12427 9331 12543 ne
tri 9331 12427 9471 12567 sw
tri 12473 12543 12497 12567 se
rect 12497 12543 12613 12567
tri 12613 12543 12637 12567 nw
rect 14566 12566 14774 14566
tri 12357 12427 12473 12543 se
tri 9331 12403 9355 12427 ne
rect 9355 12403 9471 12427
tri 6913 12287 7029 12403 se
tri 4167 12147 4307 12287 ne
tri 4307 12147 4447 12287 sw
tri 6889 12263 6913 12287 se
rect 6913 12263 7029 12287
tri 7029 12263 7169 12403 nw
tri 9355 12287 9471 12403 ne
tri 9471 12287 9611 12427 sw
tri 12333 12403 12357 12427 se
rect 12357 12403 12473 12427
tri 12473 12403 12613 12543 nw
tri 12217 12287 12333 12403 se
tri 9471 12263 9495 12287 ne
rect 9495 12263 9611 12287
tri 6773 12147 6889 12263 se
tri 4307 12007 4447 12147 ne
tri 4447 12007 4587 12147 sw
tri 6749 12123 6773 12147 se
rect 6773 12123 6889 12147
tri 6889 12123 7029 12263 nw
tri 9495 12147 9611 12263 ne
tri 9611 12147 9751 12287 sw
tri 12193 12263 12217 12287 se
rect 12217 12263 12333 12287
tri 12333 12263 12473 12403 nw
tri 12077 12147 12193 12263 se
tri 9611 12123 9635 12147 ne
rect 9635 12123 9751 12147
tri 6633 12007 6749 12123 se
tri 4447 11914 4540 12007 ne
rect 4540 11914 4587 12007
rect 1750 9914 1958 11914
tri 4540 11867 4587 11914 ne
tri 4587 11913 4681 12007 sw
tri 6609 11983 6633 12007 se
rect 6633 11983 6749 12007
tri 6749 11983 6889 12123 nw
tri 9635 12007 9751 12123 ne
tri 9751 12007 9891 12147 sw
tri 12053 12123 12077 12147 se
rect 12077 12123 12193 12147
tri 12193 12123 12333 12263 nw
tri 11937 12007 12053 12123 se
tri 9751 11983 9775 12007 ne
rect 9775 11983 9891 12007
rect 4587 11867 4611 11913
tri 4587 11843 4611 11867 ne
tri 4611 11843 4681 11913 nw
tri 6539 11913 6609 11983 se
tri 6539 11843 6609 11913 ne
tri 6609 11843 6749 11983 nw
tri 9775 11867 9891 11983 ne
tri 9891 11913 9985 12007 sw
tri 11913 11983 11937 12007 se
rect 11937 11983 12053 12007
tri 12053 11983 12193 12123 nw
rect 9891 11867 9915 11913
tri 9891 11843 9915 11867 ne
tri 9915 11843 9985 11913 nw
tri 11843 11913 11913 11983 se
tri 11843 11843 11913 11913 ne
tri 11913 11843 12053 11983 nw
tri 3887 9915 3957 9985 se
tri 3957 9915 4027 9985 sw
tri 7193 9915 7263 9985 se
tri 7263 9915 7333 9985 sw
tri 3887 9914 3888 9915 ne
rect 3888 9914 4027 9915
rect 1750 6610 1838 9914
tri 3888 9775 4027 9914 ne
tri 4027 9775 4167 9915 sw
tri 7169 9891 7193 9915 se
rect 7193 9891 7309 9915
tri 7309 9891 7333 9915 nw
tri 9191 9915 9261 9985 se
tri 9261 9915 9331 9985 sw
tri 12497 9915 12567 9985 se
tri 12567 9915 12637 9985 sw
tri 9191 9891 9215 9915 ne
rect 9215 9891 9331 9915
tri 7053 9775 7169 9891 se
tri 4027 9635 4167 9775 ne
tri 4167 9635 4307 9775 sw
tri 7029 9751 7053 9775 se
rect 7053 9751 7169 9775
tri 7169 9751 7309 9891 nw
tri 9215 9775 9331 9891 ne
tri 9331 9775 9471 9915 sw
tri 12473 9891 12497 9915 se
rect 12497 9891 12613 9915
tri 12613 9891 12637 9915 nw
tri 12357 9775 12473 9891 se
tri 9331 9751 9355 9775 ne
rect 9355 9751 9471 9775
tri 6913 9635 7029 9751 se
tri 4167 9495 4307 9635 ne
tri 4307 9495 4447 9635 sw
tri 6889 9611 6913 9635 se
rect 6913 9611 7029 9635
tri 7029 9611 7169 9751 nw
tri 9355 9635 9471 9751 ne
tri 9471 9635 9611 9775 sw
tri 12333 9751 12357 9775 se
rect 12357 9751 12473 9775
tri 12473 9751 12613 9891 nw
tri 12217 9635 12333 9751 se
tri 9471 9611 9495 9635 ne
rect 9495 9611 9611 9635
tri 6773 9495 6889 9611 se
tri 4307 9355 4447 9495 ne
tri 4447 9355 4587 9495 sw
tri 6749 9471 6773 9495 se
rect 6773 9471 6889 9495
tri 6889 9471 7029 9611 nw
tri 9495 9495 9611 9611 ne
tri 9611 9495 9751 9635 sw
tri 12193 9611 12217 9635 se
rect 12217 9611 12333 9635
tri 12333 9611 12473 9751 nw
tri 12077 9495 12193 9611 se
tri 9611 9471 9635 9495 ne
rect 9635 9471 9751 9495
tri 6633 9355 6749 9471 se
tri 4447 9215 4587 9355 ne
tri 4587 9261 4681 9355 sw
tri 6609 9331 6633 9355 se
rect 6633 9331 6749 9355
tri 6749 9331 6889 9471 nw
tri 9635 9355 9751 9471 ne
tri 9751 9355 9891 9495 sw
tri 12053 9471 12077 9495 se
rect 12077 9471 12193 9495
tri 12193 9471 12333 9611 nw
tri 11937 9355 12053 9471 se
tri 9751 9331 9775 9355 ne
rect 9775 9331 9891 9355
rect 4587 9215 4611 9261
tri 4587 9191 4611 9215 ne
tri 4611 9191 4681 9261 nw
tri 6539 9261 6609 9331 se
tri 6539 9191 6609 9261 ne
tri 6609 9191 6749 9331 nw
tri 9775 9215 9891 9331 ne
tri 9891 9261 9985 9355 sw
tri 11913 9331 11937 9355 se
rect 11937 9331 12053 9355
tri 12053 9331 12193 9471 nw
rect 9891 9215 9915 9261
tri 9891 9191 9915 9215 ne
tri 9915 9191 9985 9261 nw
tri 11843 9261 11913 9331 se
tri 11843 9191 11913 9261 ne
tri 11913 9191 12053 9331 nw
rect 14686 9262 14774 12566
tri 3887 7263 3957 7333 se
tri 3957 7263 4027 7333 sw
tri 7193 7263 7263 7333 se
tri 7263 7263 7333 7333 sw
tri 3887 7123 4027 7263 ne
tri 4027 7123 4167 7263 sw
tri 7169 7239 7193 7263 se
rect 7193 7239 7309 7263
tri 7309 7239 7333 7263 nw
tri 9191 7263 9261 7333 se
tri 9261 7263 9331 7333 sw
tri 12497 7263 12567 7333 se
tri 12567 7263 12637 7333 sw
tri 9191 7239 9215 7263 ne
rect 9215 7239 9331 7263
tri 7053 7123 7169 7239 se
tri 4027 6983 4167 7123 ne
tri 4167 6983 4307 7123 sw
tri 7029 7099 7053 7123 se
rect 7053 7099 7169 7123
tri 7169 7099 7309 7239 nw
tri 9215 7123 9331 7239 ne
tri 9331 7123 9471 7263 sw
tri 12473 7239 12497 7263 se
rect 12497 7239 12613 7263
tri 12613 7239 12637 7263 nw
rect 14566 7262 14774 9262
tri 12357 7123 12473 7239 se
tri 9331 7099 9355 7123 ne
rect 9355 7099 9471 7123
tri 6913 6983 7029 7099 se
tri 4167 6843 4307 6983 ne
tri 4307 6843 4447 6983 sw
tri 6889 6959 6913 6983 se
rect 6913 6959 7029 6983
tri 7029 6959 7169 7099 nw
tri 9355 6983 9471 7099 ne
tri 9471 6983 9611 7123 sw
tri 12333 7099 12357 7123 se
rect 12357 7099 12473 7123
tri 12473 7099 12613 7239 nw
tri 12217 6983 12333 7099 se
tri 9471 6959 9495 6983 ne
rect 9495 6959 9611 6983
tri 6773 6843 6889 6959 se
tri 4307 6703 4447 6843 ne
tri 4447 6703 4587 6843 sw
tri 6749 6819 6773 6843 se
rect 6773 6819 6889 6843
tri 6889 6819 7029 6959 nw
tri 9495 6843 9611 6959 ne
tri 9611 6843 9751 6983 sw
tri 12193 6959 12217 6983 se
rect 12217 6959 12333 6983
tri 12333 6959 12473 7099 nw
tri 12077 6843 12193 6959 se
tri 9611 6819 9635 6843 ne
rect 9635 6819 9751 6843
tri 6633 6703 6749 6819 se
tri 4447 6610 4540 6703 ne
rect 4540 6610 4587 6703
rect 1750 4610 1958 6610
tri 4540 6563 4587 6610 ne
tri 4587 6609 4681 6703 sw
tri 6609 6679 6633 6703 se
rect 6633 6679 6749 6703
tri 6749 6679 6889 6819 nw
tri 9635 6703 9751 6819 ne
tri 9751 6703 9891 6843 sw
tri 12053 6819 12077 6843 se
rect 12077 6819 12193 6843
tri 12193 6819 12333 6959 nw
tri 11937 6703 12053 6819 se
tri 9751 6679 9775 6703 ne
rect 9775 6679 9891 6703
rect 4587 6563 4611 6609
tri 4587 6539 4611 6563 ne
tri 4611 6539 4681 6609 nw
tri 6539 6609 6609 6679 se
tri 6539 6539 6609 6609 ne
tri 6609 6539 6749 6679 nw
tri 9775 6563 9891 6679 ne
tri 9891 6609 9985 6703 sw
tri 11913 6679 11937 6703 se
rect 11937 6679 12053 6703
tri 12053 6679 12193 6819 nw
rect 9891 6563 9915 6609
tri 9891 6539 9915 6563 ne
tri 9915 6539 9985 6609 nw
tri 11843 6609 11913 6679 se
tri 11843 6539 11913 6609 ne
tri 11913 6539 12053 6679 nw
tri 3887 4611 3957 4681 se
tri 3957 4611 4027 4681 sw
tri 7193 4611 7263 4681 se
tri 7263 4611 7333 4681 sw
tri 3887 4610 3888 4611 ne
rect 3888 4610 4027 4611
rect 1542 1630 1630 4542
tri 3888 4471 4027 4610 ne
tri 4027 4471 4167 4611 sw
tri 7169 4587 7193 4611 se
rect 7193 4587 7309 4611
tri 7309 4587 7333 4611 nw
tri 9191 4611 9261 4681 se
tri 9261 4611 9331 4681 sw
tri 12497 4611 12567 4681 se
tri 12567 4611 12637 4681 sw
tri 9191 4587 9215 4611 ne
rect 9215 4587 9331 4611
tri 7053 4471 7169 4587 se
tri 4027 4331 4167 4471 ne
tri 4167 4331 4307 4471 sw
tri 7029 4447 7053 4471 se
rect 7053 4447 7169 4471
tri 7169 4447 7309 4587 nw
tri 9215 4471 9331 4587 ne
tri 9331 4471 9471 4611 sw
tri 12473 4587 12497 4611 se
rect 12497 4587 12613 4611
tri 12613 4587 12637 4611 nw
tri 12357 4471 12473 4587 se
tri 9331 4447 9355 4471 ne
rect 9355 4447 9471 4471
tri 6913 4331 7029 4447 se
tri 4167 4191 4307 4331 ne
tri 4307 4191 4447 4331 sw
tri 6889 4307 6913 4331 se
rect 6913 4307 7029 4331
tri 7029 4307 7169 4447 nw
tri 9355 4331 9471 4447 ne
tri 9471 4331 9611 4471 sw
tri 12333 4447 12357 4471 se
rect 12357 4447 12473 4471
tri 12473 4447 12613 4587 nw
tri 12217 4331 12333 4447 se
tri 9471 4307 9495 4331 ne
rect 9495 4307 9611 4331
tri 6773 4191 6889 4307 se
tri 4307 4051 4447 4191 ne
tri 4447 4051 4587 4191 sw
tri 6749 4167 6773 4191 se
rect 6773 4167 6889 4191
tri 6889 4167 7029 4307 nw
tri 9495 4191 9611 4307 ne
tri 9611 4191 9751 4331 sw
tri 12193 4307 12217 4331 se
rect 12217 4307 12333 4331
tri 12333 4307 12473 4447 nw
tri 12077 4191 12193 4307 se
tri 9611 4167 9635 4191 ne
rect 9635 4167 9751 4191
tri 6633 4051 6749 4167 se
tri 4447 3911 4587 4051 ne
tri 4587 3957 4681 4051 sw
tri 6609 4027 6633 4051 se
rect 6633 4027 6749 4051
tri 6749 4027 6889 4167 nw
tri 9635 4051 9751 4167 ne
tri 9751 4051 9891 4191 sw
tri 12053 4167 12077 4191 se
rect 12077 4167 12193 4191
tri 12193 4167 12333 4307 nw
tri 11937 4051 12053 4167 se
tri 9751 4027 9775 4051 ne
rect 9775 4027 9891 4051
rect 4587 3911 4611 3957
tri 4587 3887 4611 3911 ne
tri 4611 3887 4681 3957 nw
tri 6539 3957 6609 4027 se
tri 6539 3887 6609 3957 ne
tri 6609 3887 6749 4027 nw
tri 9775 3911 9891 4027 ne
tri 9891 3957 9985 4051 sw
tri 11913 4027 11937 4051 se
rect 11937 4027 12053 4051
tri 12053 4027 12193 4167 nw
rect 9891 3911 9915 3957
tri 9891 3887 9915 3911 ne
tri 9915 3887 9985 3957 nw
tri 11843 3957 11913 4027 se
tri 11843 3887 11913 3957 ne
tri 11913 3887 12053 4027 nw
rect 14686 3958 14774 7262
rect 14566 1958 14774 3958
rect 14894 30546 14982 36415
rect 14894 28410 14910 30546
rect 14966 28410 14982 30546
rect 14894 25242 14982 28410
rect 14894 23418 14910 25242
rect 14966 23418 14982 25242
rect 14894 19938 14982 23418
rect 14894 17802 14910 19938
rect 14966 17802 14982 19938
rect 14894 14634 14982 17802
rect 14894 12810 14910 14634
rect 14966 12810 14982 14634
rect 14894 9330 14982 12810
rect 14894 7194 14910 9330
rect 14966 7194 14982 9330
rect 14894 4026 14982 7194
rect 14894 2202 14910 4026
rect 14966 2202 14982 4026
rect 14894 2180 14982 2202
rect 15860 30988 15948 34512
rect 15860 30620 15876 30988
rect 15932 30620 15948 30988
rect 15860 28336 15948 30620
rect 15860 27968 15876 28336
rect 15932 27968 15948 28336
rect 15860 25684 15948 27968
rect 15860 25316 15876 25684
rect 15932 25316 15948 25684
rect 15860 23032 15948 25316
rect 15860 22664 15876 23032
rect 15932 22664 15948 23032
rect 15860 20380 15948 22664
rect 15860 20012 15876 20380
rect 15932 20012 15948 20380
rect 15860 17728 15948 20012
rect 15860 17360 15876 17728
rect 15932 17360 15948 17728
rect 15860 15076 15948 17360
rect 15860 14708 15876 15076
rect 15932 14708 15948 15076
rect 15860 12424 15948 14708
rect 15860 12056 15876 12424
rect 15932 12056 15948 12424
rect 15860 9772 15948 12056
rect 15860 9404 15876 9772
rect 15932 9404 15948 9772
rect 15860 7120 15948 9404
rect 15860 6752 15876 7120
rect 15932 6752 15948 7120
rect 15860 4468 15948 6752
rect 15860 4100 15876 4468
rect 15932 4100 15948 4468
rect 1958 1838 3958 1958
rect 7262 1838 9262 1958
rect 12566 1838 14774 1958
rect 1958 1750 14774 1838
rect 1542 1614 12034 1630
rect 1542 1558 4542 1614
rect 6678 1558 9846 1614
rect 11982 1558 12034 1614
rect 1542 1542 12034 1558
rect 15860 664 15948 4100
rect 576 648 15948 664
rect 576 592 4100 648
rect 4468 592 6752 648
rect 7120 592 9404 648
rect 9772 592 12056 648
rect 12424 592 15948 648
rect 576 576 15948 592
use cap_mim$1  cap_mim$1_0
timestamp 1587330750
transform 1 0 12566 0 1 7262
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_1
timestamp 1587330750
transform 1 0 12566 0 1 9914
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_2
timestamp 1587330750
transform 1 0 12566 0 1 1958
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_3
timestamp 1587330750
transform 1 0 12566 0 1 4610
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_4
timestamp 1587330750
transform 1 0 9914 0 1 7262
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_5
timestamp 1587330750
transform 1 0 7262 0 1 7262
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_6
timestamp 1587330750
transform 1 0 9914 0 1 9914
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_7
timestamp 1587330750
transform 1 0 7262 0 1 9914
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_8
timestamp 1587330750
transform 1 0 9914 0 1 1958
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_9
timestamp 1587330750
transform 1 0 7262 0 1 1958
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_10
timestamp 1587330750
transform 1 0 9914 0 1 4610
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_11
timestamp 1587330750
transform 1 0 7262 0 1 4610
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_12
timestamp 1587330750
transform 1 0 4610 0 1 7262
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_13
timestamp 1587330750
transform 1 0 1958 0 1 7262
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_14
timestamp 1587330750
transform 1 0 4610 0 1 9914
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_15
timestamp 1587330750
transform 1 0 1958 0 1 9914
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_16
timestamp 1587330750
transform 1 0 4610 0 1 1958
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_17
timestamp 1587330750
transform 1 0 1958 0 1 1958
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_18
timestamp 1587330750
transform 1 0 4610 0 1 4610
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_19
timestamp 1587330750
transform 1 0 1958 0 1 4610
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_20
timestamp 1587330750
transform 1 0 12566 0 1 17870
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_21
timestamp 1587330750
transform 1 0 12566 0 1 20522
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_22
timestamp 1587330750
transform 1 0 12566 0 1 12566
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_23
timestamp 1587330750
transform 1 0 12566 0 1 15218
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_24
timestamp 1587330750
transform 1 0 9914 0 1 17870
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_25
timestamp 1587330750
transform 1 0 7262 0 1 17870
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_26
timestamp 1587330750
transform 1 0 9914 0 1 20522
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_27
timestamp 1587330750
transform 1 0 7262 0 1 20522
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_28
timestamp 1587330750
transform 1 0 9914 0 1 12566
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_29
timestamp 1587330750
transform 1 0 7262 0 1 12566
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_30
timestamp 1587330750
transform 1 0 9914 0 1 15218
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_31
timestamp 1587330750
transform 1 0 7262 0 1 15218
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_32
timestamp 1587330750
transform 1 0 4610 0 1 17870
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_33
timestamp 1587330750
transform 1 0 1958 0 1 17870
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_34
timestamp 1587330750
transform 1 0 4610 0 1 20522
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_35
timestamp 1587330750
transform 1 0 1958 0 1 20522
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_36
timestamp 1587330750
transform 1 0 4610 0 1 12566
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_37
timestamp 1587330750
transform 1 0 1958 0 1 12566
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_38
timestamp 1587330750
transform 1 0 4610 0 1 15218
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_39
timestamp 1587330750
transform 1 0 1958 0 1 15218
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_40
timestamp 1587330750
transform 1 0 12566 0 1 28478
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_41
timestamp 1587330750
transform 1 0 12566 0 1 31130
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_42
timestamp 1587330750
transform 1 0 12566 0 1 23174
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_43
timestamp 1587330750
transform 1 0 12566 0 1 25826
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_44
timestamp 1587330750
transform 1 0 9914 0 1 28478
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_45
timestamp 1587330750
transform 1 0 7262 0 1 28478
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_46
timestamp 1587330750
transform 1 0 9914 0 1 31130
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_47
timestamp 1587330750
transform 1 0 7262 0 1 31130
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_48
timestamp 1587330750
transform 1 0 9914 0 1 23174
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_49
timestamp 1587330750
transform 1 0 7262 0 1 23174
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_50
timestamp 1587330750
transform 1 0 9914 0 1 25826
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_51
timestamp 1587330750
transform 1 0 7262 0 1 25826
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_52
timestamp 1587330750
transform 1 0 4610 0 1 28478
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_53
timestamp 1587330750
transform 1 0 1958 0 1 28478
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_54
timestamp 1587330750
transform 1 0 4610 0 1 31130
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_55
timestamp 1587330750
transform 1 0 1958 0 1 31130
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_56
timestamp 1587330750
transform 1 0 4610 0 1 23174
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_57
timestamp 1587330750
transform 1 0 1958 0 1 23174
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_58
timestamp 1587330750
transform 1 0 4610 0 1 25826
box -120 -120 2120 2120
use cap_mim$1  cap_mim$1_59
timestamp 1587330750
transform 1 0 1958 0 1 25826
box -120 -120 2120 2120
use cap_mim$2  cap_mim$2_0
timestamp 1587330750
transform 1 0 120 0 1 120
box -120 -120 1120 1120
use cap_mim$2  cap_mim$2_1
timestamp 1587330750
transform 1 0 15404 0 1 120
box -120 -120 1120 1120
use cap_mim$2  cap_mim$2_2
timestamp 1587330750
transform 1 0 120 0 1 33968
box -120 -120 1120 1120
use cap_mim$2  cap_mim$2_3
timestamp 1587330750
transform 1 0 15404 0 1 33968
box -120 -120 1120 1120
use cap_mim  cap_mim_0
timestamp 1587330750
transform 0 -1 14566 1 0 120
box -120 -120 1120 2120
use cap_mim  cap_mim_1
timestamp 1587330750
transform 0 -1 11914 1 0 120
box -120 -120 1120 2120
use cap_mim  cap_mim_2
timestamp 1587330750
transform 0 -1 9262 1 0 120
box -120 -120 1120 2120
use cap_mim  cap_mim_3
timestamp 1587330750
transform 0 -1 6610 1 0 120
box -120 -120 1120 2120
use cap_mim  cap_mim_4
timestamp 1587330750
transform 0 -1 3958 1 0 120
box -120 -120 1120 2120
use cap_mim  cap_mim_5
timestamp 1587330750
transform 1 0 120 0 1 1958
box -120 -120 1120 2120
use cap_mim  cap_mim_6
timestamp 1587330750
transform 1 0 120 0 1 4610
box -120 -120 1120 2120
use cap_mim  cap_mim_7
timestamp 1587330750
transform 1 0 120 0 1 7262
box -120 -120 1120 2120
use cap_mim  cap_mim_8
timestamp 1587330750
transform 1 0 120 0 1 9914
box -120 -120 1120 2120
use cap_mim  cap_mim_9
timestamp 1587330750
transform 1 0 120 0 1 12566
box -120 -120 1120 2120
use cap_mim  cap_mim_10
timestamp 1587330750
transform 1 0 120 0 1 15218
box -120 -120 1120 2120
use cap_mim  cap_mim_11
timestamp 1587330750
transform 1 0 120 0 1 17870
box -120 -120 1120 2120
use cap_mim  cap_mim_12
timestamp 1587330750
transform 1 0 120 0 1 20522
box -120 -120 1120 2120
use cap_mim  cap_mim_13
timestamp 1587330750
transform 1 0 15404 0 1 1958
box -120 -120 1120 2120
use cap_mim  cap_mim_14
timestamp 1587330750
transform 1 0 15404 0 1 4610
box -120 -120 1120 2120
use cap_mim  cap_mim_15
timestamp 1587330750
transform 1 0 15404 0 1 7262
box -120 -120 1120 2120
use cap_mim  cap_mim_16
timestamp 1587330750
transform 1 0 15404 0 1 9914
box -120 -120 1120 2120
use cap_mim  cap_mim_17
timestamp 1587330750
transform 1 0 15404 0 1 12566
box -120 -120 1120 2120
use cap_mim  cap_mim_18
timestamp 1587330750
transform 1 0 15404 0 1 15218
box -120 -120 1120 2120
use cap_mim  cap_mim_19
timestamp 1587330750
transform 1 0 15404 0 1 17870
box -120 -120 1120 2120
use cap_mim  cap_mim_20
timestamp 1587330750
transform 1 0 15404 0 1 20522
box -120 -120 1120 2120
use cap_mim  cap_mim_21
timestamp 1587330750
transform 1 0 120 0 1 23174
box -120 -120 1120 2120
use cap_mim  cap_mim_22
timestamp 1587330750
transform 1 0 120 0 1 25826
box -120 -120 1120 2120
use cap_mim  cap_mim_23
timestamp 1587330750
transform 1 0 120 0 1 28478
box -120 -120 1120 2120
use cap_mim  cap_mim_24
timestamp 1587330750
transform 1 0 120 0 1 31130
box -120 -120 1120 2120
use cap_mim  cap_mim_25
timestamp 1587330750
transform 0 -1 14566 1 0 33968
box -120 -120 1120 2120
use cap_mim  cap_mim_26
timestamp 1587330750
transform 0 -1 11914 1 0 33968
box -120 -120 1120 2120
use cap_mim  cap_mim_27
timestamp 1587330750
transform 0 -1 9262 1 0 33968
box -120 -120 1120 2120
use cap_mim  cap_mim_28
timestamp 1587330750
transform 0 -1 6610 1 0 33968
box -120 -120 1120 2120
use cap_mim  cap_mim_29
timestamp 1587330750
transform 0 -1 3958 1 0 33968
box -120 -120 1120 2120
use cap_mim  cap_mim_30
timestamp 1587330750
transform 1 0 15404 0 1 23174
box -120 -120 1120 2120
use cap_mim  cap_mim_31
timestamp 1587330750
transform 1 0 15404 0 1 25826
box -120 -120 1120 2120
use cap_mim  cap_mim_32
timestamp 1587330750
transform 1 0 15404 0 1 28478
box -120 -120 1120 2120
use cap_mim  cap_mim_33
timestamp 1587330750
transform 1 0 15404 0 1 31130
box -120 -120 1120 2120
<< labels >>
flabel metal5 s 14942 35477 14942 35477 2 FreeSans 600 0 0 0 B2
port 1 nsew
flabel metal5 s 14713 35493 14713 35493 2 FreeSans 600 0 0 0 T2
port 2 nsew
flabel metal5 s 1768 35572 1768 35572 2 FreeSans 600 0 0 0 T1
port 3 nsew
flabel metal5 s 1564 35570 1564 35570 2 FreeSans 600 0 0 0 B1
port 4 nsew
flabel metal4 s 620 33570 620 33570 0 FreeSans 1600 0 0 0 VSS
port 5 nsew
<< properties >>
string path 49.750 59.390 46.130 63.010 
<< end >>
