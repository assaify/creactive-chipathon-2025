magic
tech gf180mcuD
magscale 1 10
timestamp 1755277289
<< nwell >>
rect -806 -1210 806 1210
<< pmos >>
rect -556 -1000 -356 1000
rect -252 -1000 -52 1000
rect 52 -1000 252 1000
rect 356 -1000 556 1000
<< pdiff >>
rect -644 987 -556 1000
rect -644 -987 -631 987
rect -585 -987 -556 987
rect -644 -1000 -556 -987
rect -356 987 -252 1000
rect -356 -987 -327 987
rect -281 -987 -252 987
rect -356 -1000 -252 -987
rect -52 987 52 1000
rect -52 -987 -23 987
rect 23 -987 52 987
rect -52 -1000 52 -987
rect 252 987 356 1000
rect 252 -987 281 987
rect 327 -987 356 987
rect 252 -1000 356 -987
rect 556 987 644 1000
rect 556 -987 585 987
rect 631 -987 644 987
rect 556 -1000 644 -987
<< pdiffc >>
rect -631 -987 -585 987
rect -327 -987 -281 987
rect -23 -987 23 987
rect 281 -987 327 987
rect 585 -987 631 987
<< nsubdiff >>
rect -782 1114 782 1186
rect -782 1070 -710 1114
rect -782 -1070 -769 1070
rect -723 -1070 -710 1070
rect 710 1070 782 1114
rect -782 -1114 -710 -1070
rect 710 -1070 723 1070
rect 769 -1070 782 1070
rect 710 -1114 782 -1070
rect -782 -1186 782 -1114
<< nsubdiffcont >>
rect -769 -1070 -723 1070
rect 723 -1070 769 1070
<< polysilicon >>
rect -556 1079 -356 1092
rect -556 1033 -543 1079
rect -369 1033 -356 1079
rect -556 1000 -356 1033
rect -252 1079 -52 1092
rect -252 1033 -239 1079
rect -65 1033 -52 1079
rect -252 1000 -52 1033
rect 52 1079 252 1092
rect 52 1033 65 1079
rect 239 1033 252 1079
rect 52 1000 252 1033
rect 356 1079 556 1092
rect 356 1033 369 1079
rect 543 1033 556 1079
rect 356 1000 556 1033
rect -556 -1033 -356 -1000
rect -556 -1079 -543 -1033
rect -369 -1079 -356 -1033
rect -556 -1092 -356 -1079
rect -252 -1033 -52 -1000
rect -252 -1079 -239 -1033
rect -65 -1079 -52 -1033
rect -252 -1092 -52 -1079
rect 52 -1033 252 -1000
rect 52 -1079 65 -1033
rect 239 -1079 252 -1033
rect 52 -1092 252 -1079
rect 356 -1033 556 -1000
rect 356 -1079 369 -1033
rect 543 -1079 556 -1033
rect 356 -1092 556 -1079
<< polycontact >>
rect -543 1033 -369 1079
rect -239 1033 -65 1079
rect 65 1033 239 1079
rect 369 1033 543 1079
rect -543 -1079 -369 -1033
rect -239 -1079 -65 -1033
rect 65 -1079 239 -1033
rect 369 -1079 543 -1033
<< metal1 >>
rect -769 1127 769 1173
rect -769 1070 -723 1127
rect -554 1033 -543 1079
rect -369 1033 -358 1079
rect -250 1033 -239 1079
rect -65 1033 -54 1079
rect 54 1033 65 1079
rect 239 1033 250 1079
rect 358 1033 369 1079
rect 543 1033 554 1079
rect 723 1070 769 1127
rect -631 987 -585 998
rect -631 -998 -585 -987
rect -327 987 -281 998
rect -327 -998 -281 -987
rect -23 987 23 998
rect -23 -998 23 -987
rect 281 987 327 998
rect 281 -998 327 -987
rect 585 987 631 998
rect 585 -998 631 -987
rect -769 -1127 -723 -1070
rect -554 -1079 -543 -1033
rect -369 -1079 -358 -1033
rect -250 -1079 -239 -1033
rect -65 -1079 -54 -1033
rect 54 -1079 65 -1033
rect 239 -1079 250 -1033
rect 358 -1079 369 -1033
rect 543 -1079 554 -1033
rect 723 -1127 769 -1070
rect -769 -1173 769 -1127
<< properties >>
string FIXED_BBOX -746 -1150 746 1150
string gencell pfet_03v3
string library gf180mcu
string parameters w 10.0 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
