* Extracted by KLayout with GF180MCU LVS runset on : 08/09/2025 19:18

.SUBCKT active_load_diff_out VDD G D3 D4
M$1 D4 D4 D4 VDD pfet_03v3 L=0.8U W=7.3U AS=3.3215P AD=3.3215P PS=12.77U
+ PD=12.77U
M$2 VDD G D4 VDD pfet_03v3 L=0.8U W=14.6U AS=3.796P AD=3.796P PS=16.68U
+ PD=16.68U
M$3 D3 G VDD VDD pfet_03v3 L=0.8U W=14.6U AS=3.796P AD=3.796P PS=16.68U
+ PD=16.68U
M$7 D3 D3 D3 VDD pfet_03v3 L=0.8U W=7.3U AS=3.3215P AD=3.3215P PS=12.77U
+ PD=12.77U
.ENDS active_load_diff_out
