magic
tech gf180mcuD
magscale 1 10
timestamp 1755276408
<< pwell >>
rect -350 -6914 350 6914
<< nmos >>
rect -100 6254 100 6704
rect -100 5572 100 6022
rect -100 4890 100 5340
rect -100 4208 100 4658
rect -100 3526 100 3976
rect -100 2844 100 3294
rect -100 2162 100 2612
rect -100 1480 100 1930
rect -100 798 100 1248
rect -100 116 100 566
rect -100 -566 100 -116
rect -100 -1248 100 -798
rect -100 -1930 100 -1480
rect -100 -2612 100 -2162
rect -100 -3294 100 -2844
rect -100 -3976 100 -3526
rect -100 -4658 100 -4208
rect -100 -5340 100 -4890
rect -100 -6022 100 -5572
rect -100 -6704 100 -6254
<< ndiff >>
rect -188 6691 -100 6704
rect -188 6267 -175 6691
rect -129 6267 -100 6691
rect -188 6254 -100 6267
rect 100 6691 188 6704
rect 100 6267 129 6691
rect 175 6267 188 6691
rect 100 6254 188 6267
rect -188 6009 -100 6022
rect -188 5585 -175 6009
rect -129 5585 -100 6009
rect -188 5572 -100 5585
rect 100 6009 188 6022
rect 100 5585 129 6009
rect 175 5585 188 6009
rect 100 5572 188 5585
rect -188 5327 -100 5340
rect -188 4903 -175 5327
rect -129 4903 -100 5327
rect -188 4890 -100 4903
rect 100 5327 188 5340
rect 100 4903 129 5327
rect 175 4903 188 5327
rect 100 4890 188 4903
rect -188 4645 -100 4658
rect -188 4221 -175 4645
rect -129 4221 -100 4645
rect -188 4208 -100 4221
rect 100 4645 188 4658
rect 100 4221 129 4645
rect 175 4221 188 4645
rect 100 4208 188 4221
rect -188 3963 -100 3976
rect -188 3539 -175 3963
rect -129 3539 -100 3963
rect -188 3526 -100 3539
rect 100 3963 188 3976
rect 100 3539 129 3963
rect 175 3539 188 3963
rect 100 3526 188 3539
rect -188 3281 -100 3294
rect -188 2857 -175 3281
rect -129 2857 -100 3281
rect -188 2844 -100 2857
rect 100 3281 188 3294
rect 100 2857 129 3281
rect 175 2857 188 3281
rect 100 2844 188 2857
rect -188 2599 -100 2612
rect -188 2175 -175 2599
rect -129 2175 -100 2599
rect -188 2162 -100 2175
rect 100 2599 188 2612
rect 100 2175 129 2599
rect 175 2175 188 2599
rect 100 2162 188 2175
rect -188 1917 -100 1930
rect -188 1493 -175 1917
rect -129 1493 -100 1917
rect -188 1480 -100 1493
rect 100 1917 188 1930
rect 100 1493 129 1917
rect 175 1493 188 1917
rect 100 1480 188 1493
rect -188 1235 -100 1248
rect -188 811 -175 1235
rect -129 811 -100 1235
rect -188 798 -100 811
rect 100 1235 188 1248
rect 100 811 129 1235
rect 175 811 188 1235
rect 100 798 188 811
rect -188 553 -100 566
rect -188 129 -175 553
rect -129 129 -100 553
rect -188 116 -100 129
rect 100 553 188 566
rect 100 129 129 553
rect 175 129 188 553
rect 100 116 188 129
rect -188 -129 -100 -116
rect -188 -553 -175 -129
rect -129 -553 -100 -129
rect -188 -566 -100 -553
rect 100 -129 188 -116
rect 100 -553 129 -129
rect 175 -553 188 -129
rect 100 -566 188 -553
rect -188 -811 -100 -798
rect -188 -1235 -175 -811
rect -129 -1235 -100 -811
rect -188 -1248 -100 -1235
rect 100 -811 188 -798
rect 100 -1235 129 -811
rect 175 -1235 188 -811
rect 100 -1248 188 -1235
rect -188 -1493 -100 -1480
rect -188 -1917 -175 -1493
rect -129 -1917 -100 -1493
rect -188 -1930 -100 -1917
rect 100 -1493 188 -1480
rect 100 -1917 129 -1493
rect 175 -1917 188 -1493
rect 100 -1930 188 -1917
rect -188 -2175 -100 -2162
rect -188 -2599 -175 -2175
rect -129 -2599 -100 -2175
rect -188 -2612 -100 -2599
rect 100 -2175 188 -2162
rect 100 -2599 129 -2175
rect 175 -2599 188 -2175
rect 100 -2612 188 -2599
rect -188 -2857 -100 -2844
rect -188 -3281 -175 -2857
rect -129 -3281 -100 -2857
rect -188 -3294 -100 -3281
rect 100 -2857 188 -2844
rect 100 -3281 129 -2857
rect 175 -3281 188 -2857
rect 100 -3294 188 -3281
rect -188 -3539 -100 -3526
rect -188 -3963 -175 -3539
rect -129 -3963 -100 -3539
rect -188 -3976 -100 -3963
rect 100 -3539 188 -3526
rect 100 -3963 129 -3539
rect 175 -3963 188 -3539
rect 100 -3976 188 -3963
rect -188 -4221 -100 -4208
rect -188 -4645 -175 -4221
rect -129 -4645 -100 -4221
rect -188 -4658 -100 -4645
rect 100 -4221 188 -4208
rect 100 -4645 129 -4221
rect 175 -4645 188 -4221
rect 100 -4658 188 -4645
rect -188 -4903 -100 -4890
rect -188 -5327 -175 -4903
rect -129 -5327 -100 -4903
rect -188 -5340 -100 -5327
rect 100 -4903 188 -4890
rect 100 -5327 129 -4903
rect 175 -5327 188 -4903
rect 100 -5340 188 -5327
rect -188 -5585 -100 -5572
rect -188 -6009 -175 -5585
rect -129 -6009 -100 -5585
rect -188 -6022 -100 -6009
rect 100 -5585 188 -5572
rect 100 -6009 129 -5585
rect 175 -6009 188 -5585
rect 100 -6022 188 -6009
rect -188 -6267 -100 -6254
rect -188 -6691 -175 -6267
rect -129 -6691 -100 -6267
rect -188 -6704 -100 -6691
rect 100 -6267 188 -6254
rect 100 -6691 129 -6267
rect 175 -6691 188 -6267
rect 100 -6704 188 -6691
<< ndiffc >>
rect -175 6267 -129 6691
rect 129 6267 175 6691
rect -175 5585 -129 6009
rect 129 5585 175 6009
rect -175 4903 -129 5327
rect 129 4903 175 5327
rect -175 4221 -129 4645
rect 129 4221 175 4645
rect -175 3539 -129 3963
rect 129 3539 175 3963
rect -175 2857 -129 3281
rect 129 2857 175 3281
rect -175 2175 -129 2599
rect 129 2175 175 2599
rect -175 1493 -129 1917
rect 129 1493 175 1917
rect -175 811 -129 1235
rect 129 811 175 1235
rect -175 129 -129 553
rect 129 129 175 553
rect -175 -553 -129 -129
rect 129 -553 175 -129
rect -175 -1235 -129 -811
rect 129 -1235 175 -811
rect -175 -1917 -129 -1493
rect 129 -1917 175 -1493
rect -175 -2599 -129 -2175
rect 129 -2599 175 -2175
rect -175 -3281 -129 -2857
rect 129 -3281 175 -2857
rect -175 -3963 -129 -3539
rect 129 -3963 175 -3539
rect -175 -4645 -129 -4221
rect 129 -4645 175 -4221
rect -175 -5327 -129 -4903
rect 129 -5327 175 -4903
rect -175 -6009 -129 -5585
rect 129 -6009 175 -5585
rect -175 -6691 -129 -6267
rect 129 -6691 175 -6267
<< psubdiff >>
rect -326 6818 326 6890
rect -326 6774 -254 6818
rect -326 -6774 -313 6774
rect -267 -6774 -254 6774
rect 254 6774 326 6818
rect -326 -6818 -254 -6774
rect 254 -6774 267 6774
rect 313 -6774 326 6774
rect 254 -6818 326 -6774
rect -326 -6890 326 -6818
<< psubdiffcont >>
rect -313 -6774 -267 6774
rect 267 -6774 313 6774
<< polysilicon >>
rect -100 6783 100 6796
rect -100 6737 -87 6783
rect 87 6737 100 6783
rect -100 6704 100 6737
rect -100 6221 100 6254
rect -100 6175 -87 6221
rect 87 6175 100 6221
rect -100 6162 100 6175
rect -100 6101 100 6114
rect -100 6055 -87 6101
rect 87 6055 100 6101
rect -100 6022 100 6055
rect -100 5539 100 5572
rect -100 5493 -87 5539
rect 87 5493 100 5539
rect -100 5480 100 5493
rect -100 5419 100 5432
rect -100 5373 -87 5419
rect 87 5373 100 5419
rect -100 5340 100 5373
rect -100 4857 100 4890
rect -100 4811 -87 4857
rect 87 4811 100 4857
rect -100 4798 100 4811
rect -100 4737 100 4750
rect -100 4691 -87 4737
rect 87 4691 100 4737
rect -100 4658 100 4691
rect -100 4175 100 4208
rect -100 4129 -87 4175
rect 87 4129 100 4175
rect -100 4116 100 4129
rect -100 4055 100 4068
rect -100 4009 -87 4055
rect 87 4009 100 4055
rect -100 3976 100 4009
rect -100 3493 100 3526
rect -100 3447 -87 3493
rect 87 3447 100 3493
rect -100 3434 100 3447
rect -100 3373 100 3386
rect -100 3327 -87 3373
rect 87 3327 100 3373
rect -100 3294 100 3327
rect -100 2811 100 2844
rect -100 2765 -87 2811
rect 87 2765 100 2811
rect -100 2752 100 2765
rect -100 2691 100 2704
rect -100 2645 -87 2691
rect 87 2645 100 2691
rect -100 2612 100 2645
rect -100 2129 100 2162
rect -100 2083 -87 2129
rect 87 2083 100 2129
rect -100 2070 100 2083
rect -100 2009 100 2022
rect -100 1963 -87 2009
rect 87 1963 100 2009
rect -100 1930 100 1963
rect -100 1447 100 1480
rect -100 1401 -87 1447
rect 87 1401 100 1447
rect -100 1388 100 1401
rect -100 1327 100 1340
rect -100 1281 -87 1327
rect 87 1281 100 1327
rect -100 1248 100 1281
rect -100 765 100 798
rect -100 719 -87 765
rect 87 719 100 765
rect -100 706 100 719
rect -100 645 100 658
rect -100 599 -87 645
rect 87 599 100 645
rect -100 566 100 599
rect -100 83 100 116
rect -100 37 -87 83
rect 87 37 100 83
rect -100 24 100 37
rect -100 -37 100 -24
rect -100 -83 -87 -37
rect 87 -83 100 -37
rect -100 -116 100 -83
rect -100 -599 100 -566
rect -100 -645 -87 -599
rect 87 -645 100 -599
rect -100 -658 100 -645
rect -100 -719 100 -706
rect -100 -765 -87 -719
rect 87 -765 100 -719
rect -100 -798 100 -765
rect -100 -1281 100 -1248
rect -100 -1327 -87 -1281
rect 87 -1327 100 -1281
rect -100 -1340 100 -1327
rect -100 -1401 100 -1388
rect -100 -1447 -87 -1401
rect 87 -1447 100 -1401
rect -100 -1480 100 -1447
rect -100 -1963 100 -1930
rect -100 -2009 -87 -1963
rect 87 -2009 100 -1963
rect -100 -2022 100 -2009
rect -100 -2083 100 -2070
rect -100 -2129 -87 -2083
rect 87 -2129 100 -2083
rect -100 -2162 100 -2129
rect -100 -2645 100 -2612
rect -100 -2691 -87 -2645
rect 87 -2691 100 -2645
rect -100 -2704 100 -2691
rect -100 -2765 100 -2752
rect -100 -2811 -87 -2765
rect 87 -2811 100 -2765
rect -100 -2844 100 -2811
rect -100 -3327 100 -3294
rect -100 -3373 -87 -3327
rect 87 -3373 100 -3327
rect -100 -3386 100 -3373
rect -100 -3447 100 -3434
rect -100 -3493 -87 -3447
rect 87 -3493 100 -3447
rect -100 -3526 100 -3493
rect -100 -4009 100 -3976
rect -100 -4055 -87 -4009
rect 87 -4055 100 -4009
rect -100 -4068 100 -4055
rect -100 -4129 100 -4116
rect -100 -4175 -87 -4129
rect 87 -4175 100 -4129
rect -100 -4208 100 -4175
rect -100 -4691 100 -4658
rect -100 -4737 -87 -4691
rect 87 -4737 100 -4691
rect -100 -4750 100 -4737
rect -100 -4811 100 -4798
rect -100 -4857 -87 -4811
rect 87 -4857 100 -4811
rect -100 -4890 100 -4857
rect -100 -5373 100 -5340
rect -100 -5419 -87 -5373
rect 87 -5419 100 -5373
rect -100 -5432 100 -5419
rect -100 -5493 100 -5480
rect -100 -5539 -87 -5493
rect 87 -5539 100 -5493
rect -100 -5572 100 -5539
rect -100 -6055 100 -6022
rect -100 -6101 -87 -6055
rect 87 -6101 100 -6055
rect -100 -6114 100 -6101
rect -100 -6175 100 -6162
rect -100 -6221 -87 -6175
rect 87 -6221 100 -6175
rect -100 -6254 100 -6221
rect -100 -6737 100 -6704
rect -100 -6783 -87 -6737
rect 87 -6783 100 -6737
rect -100 -6796 100 -6783
<< polycontact >>
rect -87 6737 87 6783
rect -87 6175 87 6221
rect -87 6055 87 6101
rect -87 5493 87 5539
rect -87 5373 87 5419
rect -87 4811 87 4857
rect -87 4691 87 4737
rect -87 4129 87 4175
rect -87 4009 87 4055
rect -87 3447 87 3493
rect -87 3327 87 3373
rect -87 2765 87 2811
rect -87 2645 87 2691
rect -87 2083 87 2129
rect -87 1963 87 2009
rect -87 1401 87 1447
rect -87 1281 87 1327
rect -87 719 87 765
rect -87 599 87 645
rect -87 37 87 83
rect -87 -83 87 -37
rect -87 -645 87 -599
rect -87 -765 87 -719
rect -87 -1327 87 -1281
rect -87 -1447 87 -1401
rect -87 -2009 87 -1963
rect -87 -2129 87 -2083
rect -87 -2691 87 -2645
rect -87 -2811 87 -2765
rect -87 -3373 87 -3327
rect -87 -3493 87 -3447
rect -87 -4055 87 -4009
rect -87 -4175 87 -4129
rect -87 -4737 87 -4691
rect -87 -4857 87 -4811
rect -87 -5419 87 -5373
rect -87 -5539 87 -5493
rect -87 -6101 87 -6055
rect -87 -6221 87 -6175
rect -87 -6783 87 -6737
<< metal1 >>
rect -313 6831 313 6877
rect -313 6774 -267 6831
rect -98 6737 -87 6783
rect 87 6737 98 6783
rect 267 6774 313 6831
rect -175 6691 -129 6702
rect -175 6256 -129 6267
rect 129 6691 175 6702
rect 129 6256 175 6267
rect -98 6175 -87 6221
rect 87 6175 98 6221
rect -98 6055 -87 6101
rect 87 6055 98 6101
rect -175 6009 -129 6020
rect -175 5574 -129 5585
rect 129 6009 175 6020
rect 129 5574 175 5585
rect -98 5493 -87 5539
rect 87 5493 98 5539
rect -98 5373 -87 5419
rect 87 5373 98 5419
rect -175 5327 -129 5338
rect -175 4892 -129 4903
rect 129 5327 175 5338
rect 129 4892 175 4903
rect -98 4811 -87 4857
rect 87 4811 98 4857
rect -98 4691 -87 4737
rect 87 4691 98 4737
rect -175 4645 -129 4656
rect -175 4210 -129 4221
rect 129 4645 175 4656
rect 129 4210 175 4221
rect -98 4129 -87 4175
rect 87 4129 98 4175
rect -98 4009 -87 4055
rect 87 4009 98 4055
rect -175 3963 -129 3974
rect -175 3528 -129 3539
rect 129 3963 175 3974
rect 129 3528 175 3539
rect -98 3447 -87 3493
rect 87 3447 98 3493
rect -98 3327 -87 3373
rect 87 3327 98 3373
rect -175 3281 -129 3292
rect -175 2846 -129 2857
rect 129 3281 175 3292
rect 129 2846 175 2857
rect -98 2765 -87 2811
rect 87 2765 98 2811
rect -98 2645 -87 2691
rect 87 2645 98 2691
rect -175 2599 -129 2610
rect -175 2164 -129 2175
rect 129 2599 175 2610
rect 129 2164 175 2175
rect -98 2083 -87 2129
rect 87 2083 98 2129
rect -98 1963 -87 2009
rect 87 1963 98 2009
rect -175 1917 -129 1928
rect -175 1482 -129 1493
rect 129 1917 175 1928
rect 129 1482 175 1493
rect -98 1401 -87 1447
rect 87 1401 98 1447
rect -98 1281 -87 1327
rect 87 1281 98 1327
rect -175 1235 -129 1246
rect -175 800 -129 811
rect 129 1235 175 1246
rect 129 800 175 811
rect -98 719 -87 765
rect 87 719 98 765
rect -98 599 -87 645
rect 87 599 98 645
rect -175 553 -129 564
rect -175 118 -129 129
rect 129 553 175 564
rect 129 118 175 129
rect -98 37 -87 83
rect 87 37 98 83
rect -98 -83 -87 -37
rect 87 -83 98 -37
rect -175 -129 -129 -118
rect -175 -564 -129 -553
rect 129 -129 175 -118
rect 129 -564 175 -553
rect -98 -645 -87 -599
rect 87 -645 98 -599
rect -98 -765 -87 -719
rect 87 -765 98 -719
rect -175 -811 -129 -800
rect -175 -1246 -129 -1235
rect 129 -811 175 -800
rect 129 -1246 175 -1235
rect -98 -1327 -87 -1281
rect 87 -1327 98 -1281
rect -98 -1447 -87 -1401
rect 87 -1447 98 -1401
rect -175 -1493 -129 -1482
rect -175 -1928 -129 -1917
rect 129 -1493 175 -1482
rect 129 -1928 175 -1917
rect -98 -2009 -87 -1963
rect 87 -2009 98 -1963
rect -98 -2129 -87 -2083
rect 87 -2129 98 -2083
rect -175 -2175 -129 -2164
rect -175 -2610 -129 -2599
rect 129 -2175 175 -2164
rect 129 -2610 175 -2599
rect -98 -2691 -87 -2645
rect 87 -2691 98 -2645
rect -98 -2811 -87 -2765
rect 87 -2811 98 -2765
rect -175 -2857 -129 -2846
rect -175 -3292 -129 -3281
rect 129 -2857 175 -2846
rect 129 -3292 175 -3281
rect -98 -3373 -87 -3327
rect 87 -3373 98 -3327
rect -98 -3493 -87 -3447
rect 87 -3493 98 -3447
rect -175 -3539 -129 -3528
rect -175 -3974 -129 -3963
rect 129 -3539 175 -3528
rect 129 -3974 175 -3963
rect -98 -4055 -87 -4009
rect 87 -4055 98 -4009
rect -98 -4175 -87 -4129
rect 87 -4175 98 -4129
rect -175 -4221 -129 -4210
rect -175 -4656 -129 -4645
rect 129 -4221 175 -4210
rect 129 -4656 175 -4645
rect -98 -4737 -87 -4691
rect 87 -4737 98 -4691
rect -98 -4857 -87 -4811
rect 87 -4857 98 -4811
rect -175 -4903 -129 -4892
rect -175 -5338 -129 -5327
rect 129 -4903 175 -4892
rect 129 -5338 175 -5327
rect -98 -5419 -87 -5373
rect 87 -5419 98 -5373
rect -98 -5539 -87 -5493
rect 87 -5539 98 -5493
rect -175 -5585 -129 -5574
rect -175 -6020 -129 -6009
rect 129 -5585 175 -5574
rect 129 -6020 175 -6009
rect -98 -6101 -87 -6055
rect 87 -6101 98 -6055
rect -98 -6221 -87 -6175
rect 87 -6221 98 -6175
rect -175 -6267 -129 -6256
rect -175 -6702 -129 -6691
rect 129 -6267 175 -6256
rect 129 -6702 175 -6691
rect -313 -6831 -267 -6774
rect -98 -6783 -87 -6737
rect 87 -6783 98 -6737
rect 267 -6831 313 -6774
rect -313 -6877 313 -6831
<< properties >>
string FIXED_BBOX -290 -6854 290 6854
string gencell nfet_03v3
string library gf180mcu
string parameters w 2.25 l 1.0 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
