* NGSPICE file created from differential_load_res.ext - technology: gf180mcuD

.subckt res_cell a_80_80# a_1208_80# VSUBS
X0 a_80_80# a_1208_80# VSUBS ppolyf_u_1k r_width=1u r_length=5u
.ends

.subckt differential_load_res D3 D4 G VSS
Xres_cell_0 VSS VSS VSS res_cell
Xres_cell_1 m1_910_360# m1_1190_1892# VSS res_cell
Xres_cell_2 G m1_1202_1688# VSS res_cell
Xres_cell_3 m1_910_360# m1_630_1892# VSS res_cell
Xres_cell_4 D3 m1_642_1688# VSS res_cell
Xres_cell_5 VSS VSS VSS res_cell
Xres_cell_6 VSS VSS VSS res_cell
Xres_cell_7 m1_1202_1688# m1_1190_3400# VSS res_cell
Xres_cell_8 m1_1190_1892# m1_1202_3196# VSS res_cell
Xres_cell_9 m1_642_1688# m1_630_3400# VSS res_cell
Xres_cell_20 m1_1190_4908# m1_1202_6212# VSS res_cell
Xres_cell_21 m1_642_4704# m1_630_6416# VSS res_cell
Xres_cell_10 m1_630_1892# m1_642_3196# VSS res_cell
Xres_cell_22 m1_630_4908# m1_642_6212# VSS res_cell
Xres_cell_23 VSS VSS VSS res_cell
Xres_cell_12 VSS VSS VSS res_cell
Xres_cell_11 VSS VSS VSS res_cell
Xres_cell_24 VSS VSS VSS res_cell
Xres_cell_13 m1_1202_3196# m1_1190_4908# VSS res_cell
Xres_cell_25 m1_1202_6212# D4 VSS res_cell
Xres_cell_14 m1_1190_3400# m1_1202_4704# VSS res_cell
Xres_cell_26 m1_1190_6416# m1_630_7784# VSS res_cell
Xres_cell_15 m1_642_3196# m1_630_4908# VSS res_cell
Xres_cell_27 m1_642_6212# G VSS res_cell
Xres_cell_16 m1_630_3400# m1_642_4704# VSS res_cell
Xres_cell_28 m1_630_6416# m1_630_7784# VSS res_cell
Xres_cell_17 VSS VSS VSS res_cell
Xres_cell_29 VSS VSS VSS res_cell
Xres_cell_18 VSS VSS VSS res_cell
Xres_cell_19 m1_1202_4704# m1_1190_6416# VSS res_cell
.ends

