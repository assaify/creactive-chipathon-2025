magic
tech gf180mcuD
magscale 1 10
timestamp 1757061271
<< error_s >>
rect -2037 -440 -2035 -430
rect -2035 -450 -2025 -440
rect -2039 -496 -2037 -494
rect -2035 -496 -2025 -486
rect -2039 -506 -2035 -496
rect -2039 -635 -2037 -506
rect -1427 -742 -1425 -598
rect -1429 -752 -1425 -742
rect -1439 -762 -1429 -752
rect -1427 -754 -1425 -752
rect -256 -742 -254 -496
rect 425 -586 427 -479
rect 425 -596 429 -586
rect 425 -598 427 -596
rect 429 -606 439 -596
rect 429 -652 439 -642
rect 427 -662 429 -652
rect 1037 -742 1039 -598
rect -256 -752 -252 -742
rect 1035 -752 1039 -742
rect -256 -754 -254 -752
rect -252 -762 -242 -752
rect 1025 -762 1035 -752
rect 1037 -754 1039 -752
rect 2208 -742 2210 -496
rect 2208 -752 2212 -742
rect 2208 -754 2210 -752
rect 2212 -762 2222 -752
rect -1439 -808 -1429 -798
rect -256 -808 -254 -806
rect -252 -808 -242 -798
rect 1025 -808 1035 -798
rect 2208 -808 2210 -806
rect 2212 -808 2222 -798
rect -1429 -818 -1427 -808
rect -256 -818 -252 -808
rect 1035 -818 1037 -808
rect 2208 -818 2212 -808
rect -256 -860 -254 -818
rect 2208 -860 2210 -818
<< metal1 >>
rect -2240 -90 2464 90
rect -2240 -1098 2464 -918
<< via1 >>
rect -2089 -635 -2037 -479
rect -1427 -754 -1375 -598
rect -306 -860 -254 -496
rect 375 -635 427 -479
rect 1037 -754 1089 -598
rect 2158 -860 2210 -496
<< metal2 >>
rect -2093 -440 -2037 -406
rect -2093 -496 -2091 -440
rect 371 -479 427 -406
rect -310 -496 -254 -484
rect -2093 -635 -2089 -496
rect -2093 -701 -2037 -635
rect -1427 -598 -1371 -585
rect -1375 -752 -1371 -598
rect -1373 -808 -1371 -752
rect -1427 -820 -1371 -808
rect -310 -752 -306 -496
rect 371 -596 375 -479
rect 2154 -496 2210 -484
rect 371 -652 373 -596
rect 1037 -598 1093 -585
rect 371 -701 427 -652
rect 1089 -752 1093 -598
rect -310 -808 -308 -752
rect 1091 -808 1093 -752
rect -310 -860 -306 -808
rect 1037 -820 1093 -808
rect 2154 -752 2158 -496
rect 2154 -808 2156 -752
rect -310 -872 -254 -860
rect 2154 -860 2158 -808
rect 2154 -872 2210 -860
<< via2 >>
rect -2091 -479 -2035 -440
rect -2091 -496 -2089 -479
rect -2089 -496 -2037 -479
rect -2037 -496 -2035 -479
rect -1429 -754 -1427 -752
rect -1427 -754 -1375 -752
rect -1375 -754 -1373 -752
rect -1429 -808 -1373 -754
rect 373 -635 375 -596
rect 375 -635 427 -596
rect 427 -635 429 -596
rect 373 -652 429 -635
rect -308 -808 -306 -752
rect -306 -808 -254 -752
rect -254 -808 -252 -752
rect 1035 -754 1037 -752
rect 1037 -754 1089 -752
rect 1089 -754 1091 -752
rect 1035 -808 1091 -754
rect 2156 -808 2158 -752
rect 2158 -808 2210 -752
rect 2210 -808 2212 -752
<< metal3 >>
rect -2241 -440 2464 -418
rect -2241 -496 -2091 -440
rect -2035 -496 2464 -440
rect -2241 -518 2464 -496
rect -2241 -596 2464 -574
rect -2241 -652 373 -596
rect 429 -652 2464 -596
rect -2241 -674 2464 -652
rect -2241 -752 -1363 -730
rect -2241 -808 -1429 -752
rect -1373 -808 -1363 -752
rect -2241 -830 -1363 -808
rect -318 -752 1101 -730
rect -318 -808 -308 -752
rect -252 -808 1035 -752
rect 1091 -808 1101 -752
rect -318 -830 1101 -808
rect 2146 -752 2464 -730
rect 2146 -808 2156 -752
rect 2212 -808 2464 -752
rect 2146 -830 2464 -808
use gf180mcu_fd_sc_mcu9t5v0__filltie  gf180mcu_fd_sc_mcu9t5v0__filltie_0
timestamp 1757061271
transform 1 0 0 0 1 -1008
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_1  gf180mcu_fd_sc_mcu9t5v0__latq_1_0
timestamp 1757061271
transform 1 0 224 0 1 -1008
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_1  gf180mcu_fd_sc_mcu9t5v0__latq_1_1
timestamp 1757061271
transform 1 0 -2240 0 1 -1008
box -86 -90 2326 1098
<< labels >>
flabel metal1 s -2238 -1096 -2238 -1096 2 FreeSans 73 0 0 0 VSSD
port 1 nsew
flabel metal1 s -2238 88 -2238 88 4 FreeSans 73 0 0 0 VDDD
port 2 nsew
flabel metal3 s -2239 -468 -2239 -468 2 FreeSans 89 0 0 0 CLK_PH1
port 3 nsew
flabel metal3 s -2239 -624 -2239 -624 2 FreeSans 89 0 0 0 CLK_PH2
port 4 nsew
flabel metal3 s -2239 -780 -2239 -780 2 FreeSans 89 0 0 0 D
port 5 nsew
flabel metal3 s 2462 -780 2462 -780 8 FreeSans 89 0 0 0 Q
port 6 nsew
<< properties >>
string path -11.205 -2.340 12.320 -2.340 
<< end >>
