magic
tech gf180mcuD
magscale 1 10
timestamp 1757694669
<< psubdiff >>
rect 36 8213 2140 8240
rect 36 8167 214 8213
rect 1994 8167 2140 8213
rect 36 8140 2140 8167
rect 36 8088 136 8140
rect 36 188 63 8088
rect 109 188 136 8088
rect 36 136 136 188
rect 2040 8088 2140 8140
rect 2040 188 2067 8088
rect 2113 188 2140 8088
rect 2040 136 2140 188
rect 36 109 2140 136
rect 36 63 214 109
rect 1994 63 2140 109
rect 36 36 2140 63
<< psubdiffcont >>
rect 214 8167 1994 8213
rect 63 188 109 8088
rect 2067 188 2113 8088
rect 214 63 1994 109
<< metal1 >>
rect 0 8213 2176 8276
rect 0 8167 214 8213
rect 1994 8167 2176 8213
rect 0 8104 2176 8167
rect 0 8088 172 8104
rect 0 188 63 8088
rect 109 7784 172 8088
rect 2004 8088 2176 8104
rect 2004 7784 2067 8088
rect 109 7708 350 7784
rect 986 7772 1190 7784
rect 986 7720 1062 7772
rect 1114 7720 1190 7772
rect 986 7708 1190 7720
rect 1826 7708 2067 7784
rect 109 6600 172 7708
rect 2004 6600 2067 7708
rect 109 6524 350 6600
rect 630 6524 706 6600
tri 706 6524 738 6556 sw
rect 1190 6524 1266 6600
tri 1266 6524 1298 6556 sw
rect 1826 6524 2067 6600
rect 109 6276 172 6524
tri 630 6416 738 6524 ne
tri 738 6416 846 6524 sw
tri 1190 6416 1298 6524 ne
tri 1298 6416 1406 6524 sw
tri 738 6308 846 6416 ne
tri 846 6352 910 6416 sw
tri 1298 6352 1362 6416 ne
rect 1362 6352 1406 6416
tri 1406 6352 1470 6416 sw
rect 846 6308 910 6352
tri 846 6276 878 6308 ne
rect 878 6276 910 6308
tri 910 6276 986 6352 sw
tri 1362 6308 1406 6352 ne
rect 1406 6308 1470 6352
rect 109 6200 350 6276
tri 878 6244 910 6276 ne
rect 910 6200 986 6276
tri 1406 6244 1470 6308 ne
tri 1470 6276 1546 6352 sw
rect 2004 6276 2067 6524
rect 1470 6200 1546 6276
rect 1826 6200 2067 6276
rect 109 5092 172 6200
rect 2004 5092 2067 6200
rect 109 5016 350 5092
rect 630 5016 706 5092
tri 706 5016 738 5048 sw
rect 1190 5016 1266 5092
tri 1266 5016 1298 5048 sw
rect 1826 5016 2067 5092
rect 109 4768 172 5016
tri 630 4908 738 5016 ne
tri 738 4908 846 5016 sw
tri 1190 4908 1298 5016 ne
tri 1298 4908 1406 5016 sw
tri 738 4800 846 4908 ne
tri 846 4844 910 4908 sw
tri 1298 4844 1362 4908 ne
rect 1362 4844 1406 4908
tri 1406 4844 1470 4908 sw
rect 846 4800 910 4844
tri 846 4768 878 4800 ne
rect 878 4768 910 4800
tri 910 4768 986 4844 sw
tri 1362 4800 1406 4844 ne
rect 1406 4800 1470 4844
rect 109 4692 350 4768
tri 878 4736 910 4768 ne
rect 910 4692 986 4768
tri 1406 4736 1470 4800 ne
tri 1470 4768 1546 4844 sw
rect 2004 4768 2067 5016
rect 1470 4692 1546 4768
rect 1826 4692 2067 4768
rect 109 3584 172 4692
rect 2004 3584 2067 4692
rect 109 3508 350 3584
rect 630 3508 706 3584
tri 706 3508 738 3540 sw
rect 1190 3508 1266 3584
tri 1266 3508 1298 3540 sw
rect 1826 3508 2067 3584
rect 109 3260 172 3508
tri 630 3400 738 3508 ne
tri 738 3400 846 3508 sw
tri 1190 3400 1298 3508 ne
tri 1298 3400 1406 3508 sw
tri 738 3292 846 3400 ne
tri 846 3336 910 3400 sw
tri 1298 3336 1362 3400 ne
rect 1362 3336 1406 3400
tri 1406 3336 1470 3400 sw
rect 846 3292 910 3336
tri 846 3260 878 3292 ne
rect 878 3260 910 3292
tri 910 3260 986 3336 sw
tri 1362 3292 1406 3336 ne
rect 1406 3292 1470 3336
rect 109 3184 350 3260
tri 878 3228 910 3260 ne
rect 910 3184 986 3260
tri 1406 3228 1470 3292 ne
tri 1470 3260 1546 3336 sw
rect 2004 3260 2067 3508
rect 1470 3184 1546 3260
rect 1826 3184 2067 3260
rect 109 2076 172 3184
rect 2004 2076 2067 3184
rect 109 2000 350 2076
rect 630 2000 706 2076
tri 706 2000 738 2032 sw
rect 1190 2000 1266 2076
tri 1266 2000 1298 2032 sw
rect 1826 2000 2067 2076
rect 109 1752 172 2000
tri 630 1892 738 2000 ne
tri 738 1892 846 2000 sw
tri 1190 1892 1298 2000 ne
tri 1298 1892 1406 2000 sw
tri 738 1784 846 1892 ne
tri 846 1828 910 1892 sw
tri 1298 1828 1362 1892 ne
rect 1362 1828 1406 1892
tri 1406 1828 1470 1892 sw
rect 846 1784 910 1828
tri 846 1752 878 1784 ne
rect 878 1752 910 1784
tri 910 1752 986 1828 sw
tri 1362 1784 1406 1828 ne
rect 1406 1784 1470 1828
rect 109 1676 350 1752
tri 878 1720 910 1752 ne
rect 910 1676 986 1752
tri 1406 1720 1470 1784 ne
tri 1470 1752 1546 1828 sw
rect 2004 1752 2067 2000
rect 1470 1676 1546 1752
rect 1826 1676 2067 1752
rect 109 568 172 1676
rect 2004 568 2067 1676
rect 109 492 350 568
rect 1826 492 2067 568
rect 109 188 172 492
rect 630 292 706 492
rect 910 424 986 492
rect 910 372 922 424
rect 974 372 986 424
rect 910 360 986 372
rect 630 240 642 292
rect 694 240 706 292
rect 630 228 706 240
rect 1190 292 1266 492
rect 1470 424 1546 492
rect 1470 372 1482 424
rect 1534 372 1546 424
rect 1470 360 1546 372
rect 1190 240 1202 292
rect 1254 240 1266 292
rect 1190 228 1266 240
rect 0 172 172 188
rect 2004 188 2067 492
rect 2113 188 2176 8088
rect 2004 172 2176 188
rect 0 109 2176 172
rect 0 63 214 109
rect 1994 63 2176 109
rect 0 0 2176 63
<< via1 >>
rect 642 7720 694 7772
rect 1062 7720 1114 7772
rect 1482 7720 1534 7772
rect 922 6536 974 6588
rect 1482 6536 1534 6588
rect 642 6212 694 6264
rect 1202 6212 1254 6264
rect 922 5028 974 5080
rect 1482 5028 1534 5080
rect 642 4704 694 4756
rect 1202 4704 1254 4756
rect 922 3520 974 3572
rect 1482 3520 1534 3572
rect 642 3196 694 3248
rect 1202 3196 1254 3248
rect 922 2012 974 2064
rect 1482 2012 1534 2064
rect 642 1688 694 1740
rect 1202 1688 1254 1740
rect 922 372 974 424
rect 642 240 694 292
rect 1482 372 1534 424
rect 1202 240 1254 292
<< metal2 >>
rect 630 7772 706 8276
rect 630 7720 642 7772
rect 694 7720 706 7772
rect 630 7708 706 7720
rect 1050 7772 1126 8276
rect 1050 7720 1062 7772
rect 1114 7720 1126 7772
rect 1050 7708 1126 7720
rect 1470 7772 1546 8276
rect 1470 7720 1482 7772
rect 1534 7720 1546 7772
rect 1470 7708 1546 7720
rect 910 6588 986 6600
tri 890 6536 910 6556 se
rect 910 6536 922 6588
rect 974 6536 986 6588
rect 1470 6588 1546 6600
tri 1450 6536 1470 6556 se
rect 1470 6536 1482 6588
rect 1534 6536 1546 6588
tri 802 6448 890 6536 se
rect 890 6524 986 6536
rect 890 6448 910 6524
tri 910 6448 986 6524 nw
tri 1362 6448 1450 6536 se
rect 1450 6524 1546 6536
rect 1450 6448 1470 6524
tri 1470 6448 1546 6524 nw
tri 694 6340 802 6448 se
tri 802 6340 910 6448 nw
tri 1254 6340 1362 6448 se
tri 1362 6340 1470 6448 nw
tri 630 6276 694 6340 se
rect 694 6276 726 6340
rect 630 6264 726 6276
tri 726 6264 802 6340 nw
tri 1190 6276 1254 6340 se
rect 1254 6276 1266 6340
rect 1190 6264 1266 6276
rect 630 6212 642 6264
rect 694 6212 706 6264
tri 706 6244 726 6264 nw
rect 630 6200 706 6212
rect 1190 6212 1202 6264
rect 1254 6212 1266 6264
tri 1266 6244 1362 6340 nw
rect 1190 6200 1266 6212
rect 910 5080 986 5092
tri 890 5028 910 5048 se
rect 910 5028 922 5080
rect 974 5028 986 5080
rect 1470 5080 1546 5092
tri 1450 5028 1470 5048 se
rect 1470 5028 1482 5080
rect 1534 5028 1546 5080
tri 802 4940 890 5028 se
rect 890 5016 986 5028
rect 890 4940 910 5016
tri 910 4940 986 5016 nw
tri 1362 4940 1450 5028 se
rect 1450 5016 1546 5028
rect 1450 4940 1470 5016
tri 1470 4940 1546 5016 nw
tri 694 4832 802 4940 se
tri 802 4832 910 4940 nw
tri 1254 4832 1362 4940 se
tri 1362 4832 1470 4940 nw
tri 630 4768 694 4832 se
rect 694 4768 726 4832
rect 630 4756 726 4768
tri 726 4756 802 4832 nw
tri 1190 4768 1254 4832 se
rect 1254 4768 1266 4832
rect 1190 4756 1266 4768
rect 630 4704 642 4756
rect 694 4704 706 4756
tri 706 4736 726 4756 nw
rect 630 4692 706 4704
rect 1190 4704 1202 4756
rect 1254 4704 1266 4756
tri 1266 4736 1362 4832 nw
rect 1190 4692 1266 4704
rect 910 3572 986 3584
tri 890 3520 910 3540 se
rect 910 3520 922 3572
rect 974 3520 986 3572
rect 1470 3572 1546 3584
tri 1450 3520 1470 3540 se
rect 1470 3520 1482 3572
rect 1534 3520 1546 3572
tri 802 3432 890 3520 se
rect 890 3508 986 3520
rect 890 3432 910 3508
tri 910 3432 986 3508 nw
tri 1362 3432 1450 3520 se
rect 1450 3508 1546 3520
rect 1450 3432 1470 3508
tri 1470 3432 1546 3508 nw
tri 694 3324 802 3432 se
tri 802 3324 910 3432 nw
tri 1254 3324 1362 3432 se
tri 1362 3324 1470 3432 nw
tri 630 3260 694 3324 se
rect 694 3260 726 3324
rect 630 3248 726 3260
tri 726 3248 802 3324 nw
tri 1190 3260 1254 3324 se
rect 1254 3260 1266 3324
rect 1190 3248 1266 3260
rect 630 3196 642 3248
rect 694 3196 706 3248
tri 706 3228 726 3248 nw
rect 630 3184 706 3196
rect 1190 3196 1202 3248
rect 1254 3196 1266 3248
tri 1266 3228 1362 3324 nw
rect 1190 3184 1266 3196
rect 910 2064 986 2076
tri 890 2012 910 2032 se
rect 910 2012 922 2064
rect 974 2012 986 2064
rect 1470 2064 1546 2076
tri 1450 2012 1470 2032 se
rect 1470 2012 1482 2064
rect 1534 2012 1546 2064
tri 802 1924 890 2012 se
rect 890 2000 986 2012
rect 890 1924 910 2000
tri 910 1924 986 2000 nw
tri 1362 1924 1450 2012 se
rect 1450 2000 1546 2012
rect 1450 1924 1470 2000
tri 1470 1924 1546 2000 nw
tri 694 1816 802 1924 se
tri 802 1816 910 1924 nw
tri 1254 1816 1362 1924 se
tri 1362 1816 1470 1924 nw
tri 630 1752 694 1816 se
rect 694 1752 726 1816
rect 630 1740 726 1752
tri 726 1740 802 1816 nw
tri 1190 1752 1254 1816 se
rect 1254 1752 1266 1816
rect 1190 1740 1266 1752
rect 630 1688 642 1740
rect 694 1688 706 1740
tri 706 1720 726 1740 nw
rect 630 1676 706 1688
rect 1190 1688 1202 1740
rect 1254 1688 1266 1740
tri 1266 1720 1362 1816 nw
rect 1190 1676 1266 1688
rect 910 424 1546 436
rect 910 372 922 424
rect 974 372 1482 424
rect 1534 372 1546 424
rect 910 360 1546 372
rect 630 292 1266 304
rect 630 240 642 292
rect 694 240 1202 292
rect 1254 240 1266 292
rect 630 228 1266 240
use resss  resss_0
timestamp 1586290328
transform 0 -1 1968 1 0 414
box 78 80 1338 280
use resss  resss_1
timestamp 1586290328
transform 0 -1 1688 1 0 414
box 78 80 1338 280
use resss  resss_2
timestamp 1586290328
transform 0 -1 1408 1 0 414
box 78 80 1338 280
use resss  resss_3
timestamp 1586290328
transform 0 -1 1128 1 0 414
box 78 80 1338 280
use resss  resss_4
timestamp 1586290328
transform 0 -1 848 1 0 414
box 78 80 1338 280
use resss  resss_5
timestamp 1586290328
transform 0 -1 568 1 0 414
box 78 80 1338 280
use resss  resss_6
timestamp 1586290328
transform 0 -1 1968 1 0 1922
box 78 80 1338 280
use resss  resss_7
timestamp 1586290328
transform 0 -1 1688 1 0 1922
box 78 80 1338 280
use resss  resss_8
timestamp 1586290328
transform 0 -1 1408 1 0 1922
box 78 80 1338 280
use resss  resss_9
timestamp 1586290328
transform 0 -1 1128 1 0 1922
box 78 80 1338 280
use resss  resss_10
timestamp 1586290328
transform 0 -1 848 1 0 1922
box 78 80 1338 280
use resss  resss_11
timestamp 1586290328
transform 0 -1 568 1 0 1922
box 78 80 1338 280
use resss  resss_12
timestamp 1586290328
transform 0 -1 1968 1 0 3430
box 78 80 1338 280
use resss  resss_13
timestamp 1586290328
transform 0 -1 1688 1 0 3430
box 78 80 1338 280
use resss  resss_14
timestamp 1586290328
transform 0 -1 1408 1 0 3430
box 78 80 1338 280
use resss  resss_15
timestamp 1586290328
transform 0 -1 1128 1 0 3430
box 78 80 1338 280
use resss  resss_16
timestamp 1586290328
transform 0 -1 848 1 0 3430
box 78 80 1338 280
use resss  resss_17
timestamp 1586290328
transform 0 -1 568 1 0 3430
box 78 80 1338 280
use resss  resss_18
timestamp 1586290328
transform 0 -1 1968 1 0 4938
box 78 80 1338 280
use resss  resss_19
timestamp 1586290328
transform 0 -1 1688 1 0 4938
box 78 80 1338 280
use resss  resss_20
timestamp 1586290328
transform 0 -1 1408 1 0 4938
box 78 80 1338 280
use resss  resss_21
timestamp 1586290328
transform 0 -1 1128 1 0 4938
box 78 80 1338 280
use resss  resss_22
timestamp 1586290328
transform 0 -1 848 1 0 4938
box 78 80 1338 280
use resss  resss_23
timestamp 1586290328
transform 0 -1 568 1 0 4938
box 78 80 1338 280
use resss  resss_24
timestamp 1586290328
transform 0 -1 1968 1 0 6446
box 78 80 1338 280
use resss  resss_25
timestamp 1586290328
transform 0 -1 1688 1 0 6446
box 78 80 1338 280
use resss  resss_26
timestamp 1586290328
transform 0 -1 1408 1 0 6446
box 78 80 1338 280
use resss  resss_27
timestamp 1586290328
transform 0 -1 1128 1 0 6446
box 78 80 1338 280
use resss  resss_28
timestamp 1586290328
transform 0 -1 848 1 0 6446
box 78 80 1338 280
use resss  resss_29
timestamp 1586290328
transform 0 -1 568 1 0 6446
box 78 80 1338 280
<< labels >>
flabel metal2 s 1067 8033 1067 8033 2 FreeSans 600 0 0 0 G
port 3 nsew
flabel metal2 s 1483 8052 1483 8052 2 FreeSans 600 0 0 0 D4
port 2 nsew
flabel metal2 s 653 8054 653 8054 2 FreeSans 600 0 0 0 D3
port 1 nsew
flabel metal1 s 74 8199 74 8199 0 FreeSans 480 0 0 0 VSS
port 4 nsew
<< properties >>
string path 5.440 38.540 5.440 41.380 
<< end >>
