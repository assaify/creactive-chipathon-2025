magic
tech gf180mcuD
timestamp 1758347661
use cap_mim$1  cap_mim$1_0
timestamp 1758347661
transform 1 0 0 0 1 0
box -12 -12 212 212
<< end >>
