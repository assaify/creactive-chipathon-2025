* Extracted by KLayout with GF180MCU LVS runset on : 05/09/2025 15:33

.SUBCKT input_pair VSS D1 S D2
M$1 D1 D1 D1 VSS nfet_03v3 L=0.8U W=7.56U AS=3.2886P AD=3.2886P PS=13.08U
+ PD=13.08U
M$2 S \$3 D1 VSS nfet_03v3 L=0.8U W=15.12U AS=3.9312P AD=3.9312P PS=17.2U
+ PD=17.2U
M$3 D2 \$4 S VSS nfet_03v3 L=0.8U W=15.12U AS=3.9312P AD=3.9312P PS=17.2U
+ PD=17.2U
M$7 D2 D2 D2 VSS nfet_03v3 L=0.8U W=7.56U AS=3.2886P AD=3.2886P PS=13.08U
+ PD=13.08U
.ENDS input_pair
