* Extracted by KLayout with GF180MCU LVS runset on : 23/08/2025 09:11

.SUBCKT inv VDD OUT VSS IN
M$1 VDD IN OUT VDD pfet_03v3 L=0.28U W=1.5U AS=0.975P AD=0.975P PS=4.3U PD=4.3U
M$2 VSS IN OUT VSS nfet_03v3 L=0.28U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
.ENDS inv
