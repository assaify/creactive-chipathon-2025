magic
tech gf180mcuD
magscale 1 10
timestamp 1757061271
<< error_s >>
rect 72 761 144 771
rect 72 498 160 761
rect 72 485 144 498
rect 144 357 160 372
rect 72 294 160 357
rect 72 250 85 294
rect 124 250 160 294
rect 36 193 160 250
rect 36 147 49 193
rect 72 147 160 193
rect 36 110 160 147
rect 36 92 144 110
rect 72 82 144 92
use gf180mcu_fd_sc_mcu9t5v0__filltie  gf180mcu_fd_sc_mcu9t5v0__filltie_0
timestamp 1757061271
transform 1 0 0 0 1 0
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_1  gf180mcu_fd_sc_mcu9t5v0__latq_1_0
timestamp 1757061271
transform 1 0 0 0 1 0
box -86 -90 2326 1098
<< end >>
