magic
tech gf180mcuD
magscale 1 10
timestamp 1755255420
<< checkpaint >>
rect -2060 -2060 5086 8112
use ppolyf_u_1k_5PYHRH  XR4
timestamp 0
transform 1 0 1513 0 1 3026
box -1573 -3086 1573 3086
<< end >>
