magic
tech gf180mcuD
magscale 1 10
timestamp 1755277289
<< pwell >>
rect -806 -685 806 685
<< nmos >>
rect -556 -475 -356 475
rect -252 -475 -52 475
rect 52 -475 252 475
rect 356 -475 556 475
<< ndiff >>
rect -644 462 -556 475
rect -644 -462 -631 462
rect -585 -462 -556 462
rect -644 -475 -556 -462
rect -356 462 -252 475
rect -356 -462 -327 462
rect -281 -462 -252 462
rect -356 -475 -252 -462
rect -52 462 52 475
rect -52 -462 -23 462
rect 23 -462 52 462
rect -52 -475 52 -462
rect 252 462 356 475
rect 252 -462 281 462
rect 327 -462 356 462
rect 252 -475 356 -462
rect 556 462 644 475
rect 556 -462 585 462
rect 631 -462 644 462
rect 556 -475 644 -462
<< ndiffc >>
rect -631 -462 -585 462
rect -327 -462 -281 462
rect -23 -462 23 462
rect 281 -462 327 462
rect 585 -462 631 462
<< psubdiff >>
rect -782 589 782 661
rect -782 545 -710 589
rect -782 -545 -769 545
rect -723 -545 -710 545
rect 710 545 782 589
rect -782 -589 -710 -545
rect 710 -545 723 545
rect 769 -545 782 545
rect 710 -589 782 -545
rect -782 -661 782 -589
<< psubdiffcont >>
rect -769 -545 -723 545
rect 723 -545 769 545
<< polysilicon >>
rect -556 554 -356 567
rect -556 508 -543 554
rect -369 508 -356 554
rect -556 475 -356 508
rect -252 554 -52 567
rect -252 508 -239 554
rect -65 508 -52 554
rect -252 475 -52 508
rect 52 554 252 567
rect 52 508 65 554
rect 239 508 252 554
rect 52 475 252 508
rect 356 554 556 567
rect 356 508 369 554
rect 543 508 556 554
rect 356 475 556 508
rect -556 -508 -356 -475
rect -556 -554 -543 -508
rect -369 -554 -356 -508
rect -556 -567 -356 -554
rect -252 -508 -52 -475
rect -252 -554 -239 -508
rect -65 -554 -52 -508
rect -252 -567 -52 -554
rect 52 -508 252 -475
rect 52 -554 65 -508
rect 239 -554 252 -508
rect 52 -567 252 -554
rect 356 -508 556 -475
rect 356 -554 369 -508
rect 543 -554 556 -508
rect 356 -567 556 -554
<< polycontact >>
rect -543 508 -369 554
rect -239 508 -65 554
rect 65 508 239 554
rect 369 508 543 554
rect -543 -554 -369 -508
rect -239 -554 -65 -508
rect 65 -554 239 -508
rect 369 -554 543 -508
<< metal1 >>
rect -769 602 769 648
rect -769 545 -723 602
rect -554 508 -543 554
rect -369 508 -358 554
rect -250 508 -239 554
rect -65 508 -54 554
rect 54 508 65 554
rect 239 508 250 554
rect 358 508 369 554
rect 543 508 554 554
rect 723 545 769 602
rect -631 462 -585 473
rect -631 -473 -585 -462
rect -327 462 -281 473
rect -327 -473 -281 -462
rect -23 462 23 473
rect -23 -473 23 -462
rect 281 462 327 473
rect 281 -473 327 -462
rect 585 462 631 473
rect 585 -473 631 -462
rect -769 -602 -723 -545
rect -554 -554 -543 -508
rect -369 -554 -358 -508
rect -250 -554 -239 -508
rect -65 -554 -54 -508
rect 54 -554 65 -508
rect 239 -554 250 -508
rect 358 -554 369 -508
rect 543 -554 554 -508
rect 723 -602 769 -545
rect -769 -648 769 -602
<< properties >>
string FIXED_BBOX -746 -625 746 625
string gencell nfet_03v3
string library gf180mcu
string parameters w 4.75 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
