magic
tech gf180mcuD
magscale 1 10
timestamp 1757670462
<< nmos >>
rect 38 0 94 800
rect 198 0 254 800
rect 358 0 414 800
rect 518 0 574 800
rect 678 0 734 800
rect 838 0 894 800
<< ndiff >>
rect -84 729 38 800
rect -84 71 -65 729
rect -19 71 38 729
rect -84 0 38 71
rect 94 729 198 800
rect 94 71 123 729
rect 169 71 198 729
rect 94 0 198 71
rect 254 729 358 800
rect 254 71 283 729
rect 329 71 358 729
rect 254 0 358 71
rect 414 729 518 800
rect 414 71 443 729
rect 489 71 518 729
rect 414 0 518 71
rect 574 729 678 800
rect 574 71 603 729
rect 649 71 678 729
rect 574 0 678 71
rect 734 729 838 800
rect 734 71 763 729
rect 809 71 838 729
rect 734 0 838 71
rect 894 729 1016 800
rect 894 71 951 729
rect 997 71 1016 729
rect 894 0 1016 71
<< ndiffc >>
rect -65 71 -19 729
rect 123 71 169 729
rect 283 71 329 729
rect 443 71 489 729
rect 603 71 649 729
rect 763 71 809 729
rect 951 71 997 729
<< psubdiff >>
rect -256 922 1188 998
rect -256 -196 -180 922
rect 1112 -196 1188 922
rect -256 -272 1188 -196
<< polysilicon >>
rect 38 800 94 860
rect 198 800 254 860
rect 358 800 414 860
rect 518 800 574 860
rect 678 800 734 860
rect 838 800 894 860
rect 38 -60 94 0
rect 198 -60 254 0
rect 358 -60 414 0
rect 518 -60 574 0
rect 678 -60 734 0
rect 838 -60 894 0
rect 30 -73 102 -60
rect 30 -119 43 -73
rect 89 -119 102 -73
rect 30 -132 102 -119
rect 190 -73 262 -60
rect 190 -119 203 -73
rect 249 -119 262 -73
rect 190 -132 262 -119
rect 350 -73 422 -60
rect 350 -119 363 -73
rect 409 -119 422 -73
rect 350 -132 422 -119
rect 510 -73 582 -60
rect 510 -119 523 -73
rect 569 -119 582 -73
rect 510 -132 582 -119
rect 670 -73 742 -60
rect 670 -119 683 -73
rect 729 -119 742 -73
rect 670 -132 742 -119
rect 830 -73 902 -60
rect 830 -119 843 -73
rect 889 -119 902 -73
rect 830 -132 902 -119
<< polycontact >>
rect 43 -119 89 -73
rect 203 -119 249 -73
rect 363 -119 409 -73
rect 523 -119 569 -73
rect 683 -119 729 -73
rect 843 -119 889 -73
<< metal1 >>
rect -80 729 -4 744
rect -80 71 -65 729
rect -19 71 -4 729
rect -80 56 -4 71
rect 108 729 184 744
rect 108 71 123 729
rect 169 71 184 729
rect 108 56 184 71
rect 268 729 344 744
rect 268 71 283 729
rect 329 71 344 729
rect 268 56 344 71
rect 428 729 504 744
rect 428 71 443 729
rect 489 71 504 729
rect 428 56 504 71
rect 588 729 664 744
rect 588 71 603 729
rect 649 71 664 729
rect 588 56 664 71
rect 748 729 824 744
rect 748 71 763 729
rect 809 71 824 729
rect 748 56 824 71
rect 936 729 1012 744
rect 936 71 951 729
rect 997 71 1012 729
rect 936 56 1012 71
rect 28 -73 104 -58
rect 28 -119 43 -73
rect 89 -119 104 -73
rect 28 -134 104 -119
rect 188 -73 264 -58
rect 188 -119 203 -73
rect 249 -119 264 -73
rect 188 -134 264 -119
rect 348 -73 424 -58
rect 348 -119 363 -73
rect 409 -119 424 -73
rect 348 -134 424 -119
rect 508 -73 584 -58
rect 508 -119 523 -73
rect 569 -119 584 -73
rect 508 -134 584 -119
rect 668 -73 744 -58
rect 668 -119 683 -73
rect 729 -119 744 -73
rect 668 -134 744 -119
rect 828 -73 904 -58
rect 828 -119 843 -73
rect 889 -119 904 -73
rect 828 -134 904 -119
<< end >>
