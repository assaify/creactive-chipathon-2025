magic
tech gf180mcuD
magscale 1 10
timestamp 1758347661
use cap_mim$1  cap_mim$1_0
timestamp 1758347661
transform 1 0 -289 0 1 1025
box -120 -120 2120 2120
<< labels >>
flabel metal5 s 1630 2922 1630 2922 2 FreeSans 600 0 0 0 A
port 1 nsew
flabel metal4 s 1438 2997 1438 2997 2 FreeSans 600 0 0 0 B
port 2 nsew
<< end >>
