magic
tech gf180mcuD
magscale 1 10
timestamp 1755277289
<< mimcap >>
rect -8690 7900 -7690 7980
rect -8690 7060 -8610 7900
rect -7770 7060 -7690 7900
rect -8690 6980 -7690 7060
rect -7076 7900 -6076 7980
rect -7076 7060 -6996 7900
rect -6156 7060 -6076 7900
rect -7076 6980 -6076 7060
rect -5462 7900 -4462 7980
rect -5462 7060 -5382 7900
rect -4542 7060 -4462 7900
rect -5462 6980 -4462 7060
rect -3848 7900 -2848 7980
rect -3848 7060 -3768 7900
rect -2928 7060 -2848 7900
rect -3848 6980 -2848 7060
rect -2234 7900 -1234 7980
rect -2234 7060 -2154 7900
rect -1314 7060 -1234 7900
rect -2234 6980 -1234 7060
rect -620 7900 380 7980
rect -620 7060 -540 7900
rect 300 7060 380 7900
rect -620 6980 380 7060
rect 994 7900 1994 7980
rect 994 7060 1074 7900
rect 1914 7060 1994 7900
rect 994 6980 1994 7060
rect 2608 7900 3608 7980
rect 2608 7060 2688 7900
rect 3528 7060 3608 7900
rect 2608 6980 3608 7060
rect 4222 7900 5222 7980
rect 4222 7060 4302 7900
rect 5142 7060 5222 7900
rect 4222 6980 5222 7060
rect 5836 7900 6836 7980
rect 5836 7060 5916 7900
rect 6756 7060 6836 7900
rect 5836 6980 6836 7060
rect 7450 7900 8450 7980
rect 7450 7060 7530 7900
rect 8370 7060 8450 7900
rect 7450 6980 8450 7060
rect -8690 6540 -7690 6620
rect -8690 5700 -8610 6540
rect -7770 5700 -7690 6540
rect -8690 5620 -7690 5700
rect -7076 6540 -6076 6620
rect -7076 5700 -6996 6540
rect -6156 5700 -6076 6540
rect -7076 5620 -6076 5700
rect -5462 6540 -4462 6620
rect -5462 5700 -5382 6540
rect -4542 5700 -4462 6540
rect -5462 5620 -4462 5700
rect -3848 6540 -2848 6620
rect -3848 5700 -3768 6540
rect -2928 5700 -2848 6540
rect -3848 5620 -2848 5700
rect -2234 6540 -1234 6620
rect -2234 5700 -2154 6540
rect -1314 5700 -1234 6540
rect -2234 5620 -1234 5700
rect -620 6540 380 6620
rect -620 5700 -540 6540
rect 300 5700 380 6540
rect -620 5620 380 5700
rect 994 6540 1994 6620
rect 994 5700 1074 6540
rect 1914 5700 1994 6540
rect 994 5620 1994 5700
rect 2608 6540 3608 6620
rect 2608 5700 2688 6540
rect 3528 5700 3608 6540
rect 2608 5620 3608 5700
rect 4222 6540 5222 6620
rect 4222 5700 4302 6540
rect 5142 5700 5222 6540
rect 4222 5620 5222 5700
rect 5836 6540 6836 6620
rect 5836 5700 5916 6540
rect 6756 5700 6836 6540
rect 5836 5620 6836 5700
rect 7450 6540 8450 6620
rect 7450 5700 7530 6540
rect 8370 5700 8450 6540
rect 7450 5620 8450 5700
rect -8690 5180 -7690 5260
rect -8690 4340 -8610 5180
rect -7770 4340 -7690 5180
rect -8690 4260 -7690 4340
rect -7076 5180 -6076 5260
rect -7076 4340 -6996 5180
rect -6156 4340 -6076 5180
rect -7076 4260 -6076 4340
rect -5462 5180 -4462 5260
rect -5462 4340 -5382 5180
rect -4542 4340 -4462 5180
rect -5462 4260 -4462 4340
rect -3848 5180 -2848 5260
rect -3848 4340 -3768 5180
rect -2928 4340 -2848 5180
rect -3848 4260 -2848 4340
rect -2234 5180 -1234 5260
rect -2234 4340 -2154 5180
rect -1314 4340 -1234 5180
rect -2234 4260 -1234 4340
rect -620 5180 380 5260
rect -620 4340 -540 5180
rect 300 4340 380 5180
rect -620 4260 380 4340
rect 994 5180 1994 5260
rect 994 4340 1074 5180
rect 1914 4340 1994 5180
rect 994 4260 1994 4340
rect 2608 5180 3608 5260
rect 2608 4340 2688 5180
rect 3528 4340 3608 5180
rect 2608 4260 3608 4340
rect 4222 5180 5222 5260
rect 4222 4340 4302 5180
rect 5142 4340 5222 5180
rect 4222 4260 5222 4340
rect 5836 5180 6836 5260
rect 5836 4340 5916 5180
rect 6756 4340 6836 5180
rect 5836 4260 6836 4340
rect 7450 5180 8450 5260
rect 7450 4340 7530 5180
rect 8370 4340 8450 5180
rect 7450 4260 8450 4340
rect -8690 3820 -7690 3900
rect -8690 2980 -8610 3820
rect -7770 2980 -7690 3820
rect -8690 2900 -7690 2980
rect -7076 3820 -6076 3900
rect -7076 2980 -6996 3820
rect -6156 2980 -6076 3820
rect -7076 2900 -6076 2980
rect -5462 3820 -4462 3900
rect -5462 2980 -5382 3820
rect -4542 2980 -4462 3820
rect -5462 2900 -4462 2980
rect -3848 3820 -2848 3900
rect -3848 2980 -3768 3820
rect -2928 2980 -2848 3820
rect -3848 2900 -2848 2980
rect -2234 3820 -1234 3900
rect -2234 2980 -2154 3820
rect -1314 2980 -1234 3820
rect -2234 2900 -1234 2980
rect -620 3820 380 3900
rect -620 2980 -540 3820
rect 300 2980 380 3820
rect -620 2900 380 2980
rect 994 3820 1994 3900
rect 994 2980 1074 3820
rect 1914 2980 1994 3820
rect 994 2900 1994 2980
rect 2608 3820 3608 3900
rect 2608 2980 2688 3820
rect 3528 2980 3608 3820
rect 2608 2900 3608 2980
rect 4222 3820 5222 3900
rect 4222 2980 4302 3820
rect 5142 2980 5222 3820
rect 4222 2900 5222 2980
rect 5836 3820 6836 3900
rect 5836 2980 5916 3820
rect 6756 2980 6836 3820
rect 5836 2900 6836 2980
rect 7450 3820 8450 3900
rect 7450 2980 7530 3820
rect 8370 2980 8450 3820
rect 7450 2900 8450 2980
rect -8690 2460 -7690 2540
rect -8690 1620 -8610 2460
rect -7770 1620 -7690 2460
rect -8690 1540 -7690 1620
rect -7076 2460 -6076 2540
rect -7076 1620 -6996 2460
rect -6156 1620 -6076 2460
rect -7076 1540 -6076 1620
rect -5462 2460 -4462 2540
rect -5462 1620 -5382 2460
rect -4542 1620 -4462 2460
rect -5462 1540 -4462 1620
rect -3848 2460 -2848 2540
rect -3848 1620 -3768 2460
rect -2928 1620 -2848 2460
rect -3848 1540 -2848 1620
rect -2234 2460 -1234 2540
rect -2234 1620 -2154 2460
rect -1314 1620 -1234 2460
rect -2234 1540 -1234 1620
rect -620 2460 380 2540
rect -620 1620 -540 2460
rect 300 1620 380 2460
rect -620 1540 380 1620
rect 994 2460 1994 2540
rect 994 1620 1074 2460
rect 1914 1620 1994 2460
rect 994 1540 1994 1620
rect 2608 2460 3608 2540
rect 2608 1620 2688 2460
rect 3528 1620 3608 2460
rect 2608 1540 3608 1620
rect 4222 2460 5222 2540
rect 4222 1620 4302 2460
rect 5142 1620 5222 2460
rect 4222 1540 5222 1620
rect 5836 2460 6836 2540
rect 5836 1620 5916 2460
rect 6756 1620 6836 2460
rect 5836 1540 6836 1620
rect 7450 2460 8450 2540
rect 7450 1620 7530 2460
rect 8370 1620 8450 2460
rect 7450 1540 8450 1620
rect -8690 1100 -7690 1180
rect -8690 260 -8610 1100
rect -7770 260 -7690 1100
rect -8690 180 -7690 260
rect -7076 1100 -6076 1180
rect -7076 260 -6996 1100
rect -6156 260 -6076 1100
rect -7076 180 -6076 260
rect -5462 1100 -4462 1180
rect -5462 260 -5382 1100
rect -4542 260 -4462 1100
rect -5462 180 -4462 260
rect -3848 1100 -2848 1180
rect -3848 260 -3768 1100
rect -2928 260 -2848 1100
rect -3848 180 -2848 260
rect -2234 1100 -1234 1180
rect -2234 260 -2154 1100
rect -1314 260 -1234 1100
rect -2234 180 -1234 260
rect -620 1100 380 1180
rect -620 260 -540 1100
rect 300 260 380 1100
rect -620 180 380 260
rect 994 1100 1994 1180
rect 994 260 1074 1100
rect 1914 260 1994 1100
rect 994 180 1994 260
rect 2608 1100 3608 1180
rect 2608 260 2688 1100
rect 3528 260 3608 1100
rect 2608 180 3608 260
rect 4222 1100 5222 1180
rect 4222 260 4302 1100
rect 5142 260 5222 1100
rect 4222 180 5222 260
rect 5836 1100 6836 1180
rect 5836 260 5916 1100
rect 6756 260 6836 1100
rect 5836 180 6836 260
rect 7450 1100 8450 1180
rect 7450 260 7530 1100
rect 8370 260 8450 1100
rect 7450 180 8450 260
rect -8690 -260 -7690 -180
rect -8690 -1100 -8610 -260
rect -7770 -1100 -7690 -260
rect -8690 -1180 -7690 -1100
rect -7076 -260 -6076 -180
rect -7076 -1100 -6996 -260
rect -6156 -1100 -6076 -260
rect -7076 -1180 -6076 -1100
rect -5462 -260 -4462 -180
rect -5462 -1100 -5382 -260
rect -4542 -1100 -4462 -260
rect -5462 -1180 -4462 -1100
rect -3848 -260 -2848 -180
rect -3848 -1100 -3768 -260
rect -2928 -1100 -2848 -260
rect -3848 -1180 -2848 -1100
rect -2234 -260 -1234 -180
rect -2234 -1100 -2154 -260
rect -1314 -1100 -1234 -260
rect -2234 -1180 -1234 -1100
rect -620 -260 380 -180
rect -620 -1100 -540 -260
rect 300 -1100 380 -260
rect -620 -1180 380 -1100
rect 994 -260 1994 -180
rect 994 -1100 1074 -260
rect 1914 -1100 1994 -260
rect 994 -1180 1994 -1100
rect 2608 -260 3608 -180
rect 2608 -1100 2688 -260
rect 3528 -1100 3608 -260
rect 2608 -1180 3608 -1100
rect 4222 -260 5222 -180
rect 4222 -1100 4302 -260
rect 5142 -1100 5222 -260
rect 4222 -1180 5222 -1100
rect 5836 -260 6836 -180
rect 5836 -1100 5916 -260
rect 6756 -1100 6836 -260
rect 5836 -1180 6836 -1100
rect 7450 -260 8450 -180
rect 7450 -1100 7530 -260
rect 8370 -1100 8450 -260
rect 7450 -1180 8450 -1100
rect -8690 -1620 -7690 -1540
rect -8690 -2460 -8610 -1620
rect -7770 -2460 -7690 -1620
rect -8690 -2540 -7690 -2460
rect -7076 -1620 -6076 -1540
rect -7076 -2460 -6996 -1620
rect -6156 -2460 -6076 -1620
rect -7076 -2540 -6076 -2460
rect -5462 -1620 -4462 -1540
rect -5462 -2460 -5382 -1620
rect -4542 -2460 -4462 -1620
rect -5462 -2540 -4462 -2460
rect -3848 -1620 -2848 -1540
rect -3848 -2460 -3768 -1620
rect -2928 -2460 -2848 -1620
rect -3848 -2540 -2848 -2460
rect -2234 -1620 -1234 -1540
rect -2234 -2460 -2154 -1620
rect -1314 -2460 -1234 -1620
rect -2234 -2540 -1234 -2460
rect -620 -1620 380 -1540
rect -620 -2460 -540 -1620
rect 300 -2460 380 -1620
rect -620 -2540 380 -2460
rect 994 -1620 1994 -1540
rect 994 -2460 1074 -1620
rect 1914 -2460 1994 -1620
rect 994 -2540 1994 -2460
rect 2608 -1620 3608 -1540
rect 2608 -2460 2688 -1620
rect 3528 -2460 3608 -1620
rect 2608 -2540 3608 -2460
rect 4222 -1620 5222 -1540
rect 4222 -2460 4302 -1620
rect 5142 -2460 5222 -1620
rect 4222 -2540 5222 -2460
rect 5836 -1620 6836 -1540
rect 5836 -2460 5916 -1620
rect 6756 -2460 6836 -1620
rect 5836 -2540 6836 -2460
rect 7450 -1620 8450 -1540
rect 7450 -2460 7530 -1620
rect 8370 -2460 8450 -1620
rect 7450 -2540 8450 -2460
rect -8690 -2980 -7690 -2900
rect -8690 -3820 -8610 -2980
rect -7770 -3820 -7690 -2980
rect -8690 -3900 -7690 -3820
rect -7076 -2980 -6076 -2900
rect -7076 -3820 -6996 -2980
rect -6156 -3820 -6076 -2980
rect -7076 -3900 -6076 -3820
rect -5462 -2980 -4462 -2900
rect -5462 -3820 -5382 -2980
rect -4542 -3820 -4462 -2980
rect -5462 -3900 -4462 -3820
rect -3848 -2980 -2848 -2900
rect -3848 -3820 -3768 -2980
rect -2928 -3820 -2848 -2980
rect -3848 -3900 -2848 -3820
rect -2234 -2980 -1234 -2900
rect -2234 -3820 -2154 -2980
rect -1314 -3820 -1234 -2980
rect -2234 -3900 -1234 -3820
rect -620 -2980 380 -2900
rect -620 -3820 -540 -2980
rect 300 -3820 380 -2980
rect -620 -3900 380 -3820
rect 994 -2980 1994 -2900
rect 994 -3820 1074 -2980
rect 1914 -3820 1994 -2980
rect 994 -3900 1994 -3820
rect 2608 -2980 3608 -2900
rect 2608 -3820 2688 -2980
rect 3528 -3820 3608 -2980
rect 2608 -3900 3608 -3820
rect 4222 -2980 5222 -2900
rect 4222 -3820 4302 -2980
rect 5142 -3820 5222 -2980
rect 4222 -3900 5222 -3820
rect 5836 -2980 6836 -2900
rect 5836 -3820 5916 -2980
rect 6756 -3820 6836 -2980
rect 5836 -3900 6836 -3820
rect 7450 -2980 8450 -2900
rect 7450 -3820 7530 -2980
rect 8370 -3820 8450 -2980
rect 7450 -3900 8450 -3820
rect -8690 -4340 -7690 -4260
rect -8690 -5180 -8610 -4340
rect -7770 -5180 -7690 -4340
rect -8690 -5260 -7690 -5180
rect -7076 -4340 -6076 -4260
rect -7076 -5180 -6996 -4340
rect -6156 -5180 -6076 -4340
rect -7076 -5260 -6076 -5180
rect -5462 -4340 -4462 -4260
rect -5462 -5180 -5382 -4340
rect -4542 -5180 -4462 -4340
rect -5462 -5260 -4462 -5180
rect -3848 -4340 -2848 -4260
rect -3848 -5180 -3768 -4340
rect -2928 -5180 -2848 -4340
rect -3848 -5260 -2848 -5180
rect -2234 -4340 -1234 -4260
rect -2234 -5180 -2154 -4340
rect -1314 -5180 -1234 -4340
rect -2234 -5260 -1234 -5180
rect -620 -4340 380 -4260
rect -620 -5180 -540 -4340
rect 300 -5180 380 -4340
rect -620 -5260 380 -5180
rect 994 -4340 1994 -4260
rect 994 -5180 1074 -4340
rect 1914 -5180 1994 -4340
rect 994 -5260 1994 -5180
rect 2608 -4340 3608 -4260
rect 2608 -5180 2688 -4340
rect 3528 -5180 3608 -4340
rect 2608 -5260 3608 -5180
rect 4222 -4340 5222 -4260
rect 4222 -5180 4302 -4340
rect 5142 -5180 5222 -4340
rect 4222 -5260 5222 -5180
rect 5836 -4340 6836 -4260
rect 5836 -5180 5916 -4340
rect 6756 -5180 6836 -4340
rect 5836 -5260 6836 -5180
rect 7450 -4340 8450 -4260
rect 7450 -5180 7530 -4340
rect 8370 -5180 8450 -4340
rect 7450 -5260 8450 -5180
rect -8690 -5700 -7690 -5620
rect -8690 -6540 -8610 -5700
rect -7770 -6540 -7690 -5700
rect -8690 -6620 -7690 -6540
rect -7076 -5700 -6076 -5620
rect -7076 -6540 -6996 -5700
rect -6156 -6540 -6076 -5700
rect -7076 -6620 -6076 -6540
rect -5462 -5700 -4462 -5620
rect -5462 -6540 -5382 -5700
rect -4542 -6540 -4462 -5700
rect -5462 -6620 -4462 -6540
rect -3848 -5700 -2848 -5620
rect -3848 -6540 -3768 -5700
rect -2928 -6540 -2848 -5700
rect -3848 -6620 -2848 -6540
rect -2234 -5700 -1234 -5620
rect -2234 -6540 -2154 -5700
rect -1314 -6540 -1234 -5700
rect -2234 -6620 -1234 -6540
rect -620 -5700 380 -5620
rect -620 -6540 -540 -5700
rect 300 -6540 380 -5700
rect -620 -6620 380 -6540
rect 994 -5700 1994 -5620
rect 994 -6540 1074 -5700
rect 1914 -6540 1994 -5700
rect 994 -6620 1994 -6540
rect 2608 -5700 3608 -5620
rect 2608 -6540 2688 -5700
rect 3528 -6540 3608 -5700
rect 2608 -6620 3608 -6540
rect 4222 -5700 5222 -5620
rect 4222 -6540 4302 -5700
rect 5142 -6540 5222 -5700
rect 4222 -6620 5222 -6540
rect 5836 -5700 6836 -5620
rect 5836 -6540 5916 -5700
rect 6756 -6540 6836 -5700
rect 5836 -6620 6836 -6540
rect 7450 -5700 8450 -5620
rect 7450 -6540 7530 -5700
rect 8370 -6540 8450 -5700
rect 7450 -6620 8450 -6540
rect -8690 -7060 -7690 -6980
rect -8690 -7900 -8610 -7060
rect -7770 -7900 -7690 -7060
rect -8690 -7980 -7690 -7900
rect -7076 -7060 -6076 -6980
rect -7076 -7900 -6996 -7060
rect -6156 -7900 -6076 -7060
rect -7076 -7980 -6076 -7900
rect -5462 -7060 -4462 -6980
rect -5462 -7900 -5382 -7060
rect -4542 -7900 -4462 -7060
rect -5462 -7980 -4462 -7900
rect -3848 -7060 -2848 -6980
rect -3848 -7900 -3768 -7060
rect -2928 -7900 -2848 -7060
rect -3848 -7980 -2848 -7900
rect -2234 -7060 -1234 -6980
rect -2234 -7900 -2154 -7060
rect -1314 -7900 -1234 -7060
rect -2234 -7980 -1234 -7900
rect -620 -7060 380 -6980
rect -620 -7900 -540 -7060
rect 300 -7900 380 -7060
rect -620 -7980 380 -7900
rect 994 -7060 1994 -6980
rect 994 -7900 1074 -7060
rect 1914 -7900 1994 -7060
rect 994 -7980 1994 -7900
rect 2608 -7060 3608 -6980
rect 2608 -7900 2688 -7060
rect 3528 -7900 3608 -7060
rect 2608 -7980 3608 -7900
rect 4222 -7060 5222 -6980
rect 4222 -7900 4302 -7060
rect 5142 -7900 5222 -7060
rect 4222 -7980 5222 -7900
rect 5836 -7060 6836 -6980
rect 5836 -7900 5916 -7060
rect 6756 -7900 6836 -7060
rect 5836 -7980 6836 -7900
rect 7450 -7060 8450 -6980
rect 7450 -7900 7530 -7060
rect 8370 -7900 8450 -7060
rect 7450 -7980 8450 -7900
<< mimcapcontact >>
rect -8610 7060 -7770 7900
rect -6996 7060 -6156 7900
rect -5382 7060 -4542 7900
rect -3768 7060 -2928 7900
rect -2154 7060 -1314 7900
rect -540 7060 300 7900
rect 1074 7060 1914 7900
rect 2688 7060 3528 7900
rect 4302 7060 5142 7900
rect 5916 7060 6756 7900
rect 7530 7060 8370 7900
rect -8610 5700 -7770 6540
rect -6996 5700 -6156 6540
rect -5382 5700 -4542 6540
rect -3768 5700 -2928 6540
rect -2154 5700 -1314 6540
rect -540 5700 300 6540
rect 1074 5700 1914 6540
rect 2688 5700 3528 6540
rect 4302 5700 5142 6540
rect 5916 5700 6756 6540
rect 7530 5700 8370 6540
rect -8610 4340 -7770 5180
rect -6996 4340 -6156 5180
rect -5382 4340 -4542 5180
rect -3768 4340 -2928 5180
rect -2154 4340 -1314 5180
rect -540 4340 300 5180
rect 1074 4340 1914 5180
rect 2688 4340 3528 5180
rect 4302 4340 5142 5180
rect 5916 4340 6756 5180
rect 7530 4340 8370 5180
rect -8610 2980 -7770 3820
rect -6996 2980 -6156 3820
rect -5382 2980 -4542 3820
rect -3768 2980 -2928 3820
rect -2154 2980 -1314 3820
rect -540 2980 300 3820
rect 1074 2980 1914 3820
rect 2688 2980 3528 3820
rect 4302 2980 5142 3820
rect 5916 2980 6756 3820
rect 7530 2980 8370 3820
rect -8610 1620 -7770 2460
rect -6996 1620 -6156 2460
rect -5382 1620 -4542 2460
rect -3768 1620 -2928 2460
rect -2154 1620 -1314 2460
rect -540 1620 300 2460
rect 1074 1620 1914 2460
rect 2688 1620 3528 2460
rect 4302 1620 5142 2460
rect 5916 1620 6756 2460
rect 7530 1620 8370 2460
rect -8610 260 -7770 1100
rect -6996 260 -6156 1100
rect -5382 260 -4542 1100
rect -3768 260 -2928 1100
rect -2154 260 -1314 1100
rect -540 260 300 1100
rect 1074 260 1914 1100
rect 2688 260 3528 1100
rect 4302 260 5142 1100
rect 5916 260 6756 1100
rect 7530 260 8370 1100
rect -8610 -1100 -7770 -260
rect -6996 -1100 -6156 -260
rect -5382 -1100 -4542 -260
rect -3768 -1100 -2928 -260
rect -2154 -1100 -1314 -260
rect -540 -1100 300 -260
rect 1074 -1100 1914 -260
rect 2688 -1100 3528 -260
rect 4302 -1100 5142 -260
rect 5916 -1100 6756 -260
rect 7530 -1100 8370 -260
rect -8610 -2460 -7770 -1620
rect -6996 -2460 -6156 -1620
rect -5382 -2460 -4542 -1620
rect -3768 -2460 -2928 -1620
rect -2154 -2460 -1314 -1620
rect -540 -2460 300 -1620
rect 1074 -2460 1914 -1620
rect 2688 -2460 3528 -1620
rect 4302 -2460 5142 -1620
rect 5916 -2460 6756 -1620
rect 7530 -2460 8370 -1620
rect -8610 -3820 -7770 -2980
rect -6996 -3820 -6156 -2980
rect -5382 -3820 -4542 -2980
rect -3768 -3820 -2928 -2980
rect -2154 -3820 -1314 -2980
rect -540 -3820 300 -2980
rect 1074 -3820 1914 -2980
rect 2688 -3820 3528 -2980
rect 4302 -3820 5142 -2980
rect 5916 -3820 6756 -2980
rect 7530 -3820 8370 -2980
rect -8610 -5180 -7770 -4340
rect -6996 -5180 -6156 -4340
rect -5382 -5180 -4542 -4340
rect -3768 -5180 -2928 -4340
rect -2154 -5180 -1314 -4340
rect -540 -5180 300 -4340
rect 1074 -5180 1914 -4340
rect 2688 -5180 3528 -4340
rect 4302 -5180 5142 -4340
rect 5916 -5180 6756 -4340
rect 7530 -5180 8370 -4340
rect -8610 -6540 -7770 -5700
rect -6996 -6540 -6156 -5700
rect -5382 -6540 -4542 -5700
rect -3768 -6540 -2928 -5700
rect -2154 -6540 -1314 -5700
rect -540 -6540 300 -5700
rect 1074 -6540 1914 -5700
rect 2688 -6540 3528 -5700
rect 4302 -6540 5142 -5700
rect 5916 -6540 6756 -5700
rect 7530 -6540 8370 -5700
rect -8610 -7900 -7770 -7060
rect -6996 -7900 -6156 -7060
rect -5382 -7900 -4542 -7060
rect -3768 -7900 -2928 -7060
rect -2154 -7900 -1314 -7060
rect -540 -7900 300 -7060
rect 1074 -7900 1914 -7060
rect 2688 -7900 3528 -7060
rect 4302 -7900 5142 -7060
rect 5916 -7900 6756 -7060
rect 7530 -7900 8370 -7060
<< metal4 >>
rect -8810 8033 -7330 8100
rect -8810 7980 -7480 8033
rect -8810 6980 -8690 7980
rect -7690 6980 -7480 7980
rect -8810 6927 -7480 6980
rect -7392 6927 -7330 8033
rect -8810 6860 -7330 6927
rect -7196 8033 -5716 8100
rect -7196 7980 -5866 8033
rect -7196 6980 -7076 7980
rect -6076 6980 -5866 7980
rect -7196 6927 -5866 6980
rect -5778 6927 -5716 8033
rect -7196 6860 -5716 6927
rect -5582 8033 -4102 8100
rect -5582 7980 -4252 8033
rect -5582 6980 -5462 7980
rect -4462 6980 -4252 7980
rect -5582 6927 -4252 6980
rect -4164 6927 -4102 8033
rect -5582 6860 -4102 6927
rect -3968 8033 -2488 8100
rect -3968 7980 -2638 8033
rect -3968 6980 -3848 7980
rect -2848 6980 -2638 7980
rect -3968 6927 -2638 6980
rect -2550 6927 -2488 8033
rect -3968 6860 -2488 6927
rect -2354 8033 -874 8100
rect -2354 7980 -1024 8033
rect -2354 6980 -2234 7980
rect -1234 6980 -1024 7980
rect -2354 6927 -1024 6980
rect -936 6927 -874 8033
rect -2354 6860 -874 6927
rect -740 8033 740 8100
rect -740 7980 590 8033
rect -740 6980 -620 7980
rect 380 6980 590 7980
rect -740 6927 590 6980
rect 678 6927 740 8033
rect -740 6860 740 6927
rect 874 8033 2354 8100
rect 874 7980 2204 8033
rect 874 6980 994 7980
rect 1994 6980 2204 7980
rect 874 6927 2204 6980
rect 2292 6927 2354 8033
rect 874 6860 2354 6927
rect 2488 8033 3968 8100
rect 2488 7980 3818 8033
rect 2488 6980 2608 7980
rect 3608 6980 3818 7980
rect 2488 6927 3818 6980
rect 3906 6927 3968 8033
rect 2488 6860 3968 6927
rect 4102 8033 5582 8100
rect 4102 7980 5432 8033
rect 4102 6980 4222 7980
rect 5222 6980 5432 7980
rect 4102 6927 5432 6980
rect 5520 6927 5582 8033
rect 4102 6860 5582 6927
rect 5716 8033 7196 8100
rect 5716 7980 7046 8033
rect 5716 6980 5836 7980
rect 6836 6980 7046 7980
rect 5716 6927 7046 6980
rect 7134 6927 7196 8033
rect 5716 6860 7196 6927
rect 7330 8033 8810 8100
rect 7330 7980 8660 8033
rect 7330 6980 7450 7980
rect 8450 6980 8660 7980
rect 7330 6927 8660 6980
rect 8748 6927 8810 8033
rect 7330 6860 8810 6927
rect -8810 6673 -7330 6740
rect -8810 6620 -7480 6673
rect -8810 5620 -8690 6620
rect -7690 5620 -7480 6620
rect -8810 5567 -7480 5620
rect -7392 5567 -7330 6673
rect -8810 5500 -7330 5567
rect -7196 6673 -5716 6740
rect -7196 6620 -5866 6673
rect -7196 5620 -7076 6620
rect -6076 5620 -5866 6620
rect -7196 5567 -5866 5620
rect -5778 5567 -5716 6673
rect -7196 5500 -5716 5567
rect -5582 6673 -4102 6740
rect -5582 6620 -4252 6673
rect -5582 5620 -5462 6620
rect -4462 5620 -4252 6620
rect -5582 5567 -4252 5620
rect -4164 5567 -4102 6673
rect -5582 5500 -4102 5567
rect -3968 6673 -2488 6740
rect -3968 6620 -2638 6673
rect -3968 5620 -3848 6620
rect -2848 5620 -2638 6620
rect -3968 5567 -2638 5620
rect -2550 5567 -2488 6673
rect -3968 5500 -2488 5567
rect -2354 6673 -874 6740
rect -2354 6620 -1024 6673
rect -2354 5620 -2234 6620
rect -1234 5620 -1024 6620
rect -2354 5567 -1024 5620
rect -936 5567 -874 6673
rect -2354 5500 -874 5567
rect -740 6673 740 6740
rect -740 6620 590 6673
rect -740 5620 -620 6620
rect 380 5620 590 6620
rect -740 5567 590 5620
rect 678 5567 740 6673
rect -740 5500 740 5567
rect 874 6673 2354 6740
rect 874 6620 2204 6673
rect 874 5620 994 6620
rect 1994 5620 2204 6620
rect 874 5567 2204 5620
rect 2292 5567 2354 6673
rect 874 5500 2354 5567
rect 2488 6673 3968 6740
rect 2488 6620 3818 6673
rect 2488 5620 2608 6620
rect 3608 5620 3818 6620
rect 2488 5567 3818 5620
rect 3906 5567 3968 6673
rect 2488 5500 3968 5567
rect 4102 6673 5582 6740
rect 4102 6620 5432 6673
rect 4102 5620 4222 6620
rect 5222 5620 5432 6620
rect 4102 5567 5432 5620
rect 5520 5567 5582 6673
rect 4102 5500 5582 5567
rect 5716 6673 7196 6740
rect 5716 6620 7046 6673
rect 5716 5620 5836 6620
rect 6836 5620 7046 6620
rect 5716 5567 7046 5620
rect 7134 5567 7196 6673
rect 5716 5500 7196 5567
rect 7330 6673 8810 6740
rect 7330 6620 8660 6673
rect 7330 5620 7450 6620
rect 8450 5620 8660 6620
rect 7330 5567 8660 5620
rect 8748 5567 8810 6673
rect 7330 5500 8810 5567
rect -8810 5313 -7330 5380
rect -8810 5260 -7480 5313
rect -8810 4260 -8690 5260
rect -7690 4260 -7480 5260
rect -8810 4207 -7480 4260
rect -7392 4207 -7330 5313
rect -8810 4140 -7330 4207
rect -7196 5313 -5716 5380
rect -7196 5260 -5866 5313
rect -7196 4260 -7076 5260
rect -6076 4260 -5866 5260
rect -7196 4207 -5866 4260
rect -5778 4207 -5716 5313
rect -7196 4140 -5716 4207
rect -5582 5313 -4102 5380
rect -5582 5260 -4252 5313
rect -5582 4260 -5462 5260
rect -4462 4260 -4252 5260
rect -5582 4207 -4252 4260
rect -4164 4207 -4102 5313
rect -5582 4140 -4102 4207
rect -3968 5313 -2488 5380
rect -3968 5260 -2638 5313
rect -3968 4260 -3848 5260
rect -2848 4260 -2638 5260
rect -3968 4207 -2638 4260
rect -2550 4207 -2488 5313
rect -3968 4140 -2488 4207
rect -2354 5313 -874 5380
rect -2354 5260 -1024 5313
rect -2354 4260 -2234 5260
rect -1234 4260 -1024 5260
rect -2354 4207 -1024 4260
rect -936 4207 -874 5313
rect -2354 4140 -874 4207
rect -740 5313 740 5380
rect -740 5260 590 5313
rect -740 4260 -620 5260
rect 380 4260 590 5260
rect -740 4207 590 4260
rect 678 4207 740 5313
rect -740 4140 740 4207
rect 874 5313 2354 5380
rect 874 5260 2204 5313
rect 874 4260 994 5260
rect 1994 4260 2204 5260
rect 874 4207 2204 4260
rect 2292 4207 2354 5313
rect 874 4140 2354 4207
rect 2488 5313 3968 5380
rect 2488 5260 3818 5313
rect 2488 4260 2608 5260
rect 3608 4260 3818 5260
rect 2488 4207 3818 4260
rect 3906 4207 3968 5313
rect 2488 4140 3968 4207
rect 4102 5313 5582 5380
rect 4102 5260 5432 5313
rect 4102 4260 4222 5260
rect 5222 4260 5432 5260
rect 4102 4207 5432 4260
rect 5520 4207 5582 5313
rect 4102 4140 5582 4207
rect 5716 5313 7196 5380
rect 5716 5260 7046 5313
rect 5716 4260 5836 5260
rect 6836 4260 7046 5260
rect 5716 4207 7046 4260
rect 7134 4207 7196 5313
rect 5716 4140 7196 4207
rect 7330 5313 8810 5380
rect 7330 5260 8660 5313
rect 7330 4260 7450 5260
rect 8450 4260 8660 5260
rect 7330 4207 8660 4260
rect 8748 4207 8810 5313
rect 7330 4140 8810 4207
rect -8810 3953 -7330 4020
rect -8810 3900 -7480 3953
rect -8810 2900 -8690 3900
rect -7690 2900 -7480 3900
rect -8810 2847 -7480 2900
rect -7392 2847 -7330 3953
rect -8810 2780 -7330 2847
rect -7196 3953 -5716 4020
rect -7196 3900 -5866 3953
rect -7196 2900 -7076 3900
rect -6076 2900 -5866 3900
rect -7196 2847 -5866 2900
rect -5778 2847 -5716 3953
rect -7196 2780 -5716 2847
rect -5582 3953 -4102 4020
rect -5582 3900 -4252 3953
rect -5582 2900 -5462 3900
rect -4462 2900 -4252 3900
rect -5582 2847 -4252 2900
rect -4164 2847 -4102 3953
rect -5582 2780 -4102 2847
rect -3968 3953 -2488 4020
rect -3968 3900 -2638 3953
rect -3968 2900 -3848 3900
rect -2848 2900 -2638 3900
rect -3968 2847 -2638 2900
rect -2550 2847 -2488 3953
rect -3968 2780 -2488 2847
rect -2354 3953 -874 4020
rect -2354 3900 -1024 3953
rect -2354 2900 -2234 3900
rect -1234 2900 -1024 3900
rect -2354 2847 -1024 2900
rect -936 2847 -874 3953
rect -2354 2780 -874 2847
rect -740 3953 740 4020
rect -740 3900 590 3953
rect -740 2900 -620 3900
rect 380 2900 590 3900
rect -740 2847 590 2900
rect 678 2847 740 3953
rect -740 2780 740 2847
rect 874 3953 2354 4020
rect 874 3900 2204 3953
rect 874 2900 994 3900
rect 1994 2900 2204 3900
rect 874 2847 2204 2900
rect 2292 2847 2354 3953
rect 874 2780 2354 2847
rect 2488 3953 3968 4020
rect 2488 3900 3818 3953
rect 2488 2900 2608 3900
rect 3608 2900 3818 3900
rect 2488 2847 3818 2900
rect 3906 2847 3968 3953
rect 2488 2780 3968 2847
rect 4102 3953 5582 4020
rect 4102 3900 5432 3953
rect 4102 2900 4222 3900
rect 5222 2900 5432 3900
rect 4102 2847 5432 2900
rect 5520 2847 5582 3953
rect 4102 2780 5582 2847
rect 5716 3953 7196 4020
rect 5716 3900 7046 3953
rect 5716 2900 5836 3900
rect 6836 2900 7046 3900
rect 5716 2847 7046 2900
rect 7134 2847 7196 3953
rect 5716 2780 7196 2847
rect 7330 3953 8810 4020
rect 7330 3900 8660 3953
rect 7330 2900 7450 3900
rect 8450 2900 8660 3900
rect 7330 2847 8660 2900
rect 8748 2847 8810 3953
rect 7330 2780 8810 2847
rect -8810 2593 -7330 2660
rect -8810 2540 -7480 2593
rect -8810 1540 -8690 2540
rect -7690 1540 -7480 2540
rect -8810 1487 -7480 1540
rect -7392 1487 -7330 2593
rect -8810 1420 -7330 1487
rect -7196 2593 -5716 2660
rect -7196 2540 -5866 2593
rect -7196 1540 -7076 2540
rect -6076 1540 -5866 2540
rect -7196 1487 -5866 1540
rect -5778 1487 -5716 2593
rect -7196 1420 -5716 1487
rect -5582 2593 -4102 2660
rect -5582 2540 -4252 2593
rect -5582 1540 -5462 2540
rect -4462 1540 -4252 2540
rect -5582 1487 -4252 1540
rect -4164 1487 -4102 2593
rect -5582 1420 -4102 1487
rect -3968 2593 -2488 2660
rect -3968 2540 -2638 2593
rect -3968 1540 -3848 2540
rect -2848 1540 -2638 2540
rect -3968 1487 -2638 1540
rect -2550 1487 -2488 2593
rect -3968 1420 -2488 1487
rect -2354 2593 -874 2660
rect -2354 2540 -1024 2593
rect -2354 1540 -2234 2540
rect -1234 1540 -1024 2540
rect -2354 1487 -1024 1540
rect -936 1487 -874 2593
rect -2354 1420 -874 1487
rect -740 2593 740 2660
rect -740 2540 590 2593
rect -740 1540 -620 2540
rect 380 1540 590 2540
rect -740 1487 590 1540
rect 678 1487 740 2593
rect -740 1420 740 1487
rect 874 2593 2354 2660
rect 874 2540 2204 2593
rect 874 1540 994 2540
rect 1994 1540 2204 2540
rect 874 1487 2204 1540
rect 2292 1487 2354 2593
rect 874 1420 2354 1487
rect 2488 2593 3968 2660
rect 2488 2540 3818 2593
rect 2488 1540 2608 2540
rect 3608 1540 3818 2540
rect 2488 1487 3818 1540
rect 3906 1487 3968 2593
rect 2488 1420 3968 1487
rect 4102 2593 5582 2660
rect 4102 2540 5432 2593
rect 4102 1540 4222 2540
rect 5222 1540 5432 2540
rect 4102 1487 5432 1540
rect 5520 1487 5582 2593
rect 4102 1420 5582 1487
rect 5716 2593 7196 2660
rect 5716 2540 7046 2593
rect 5716 1540 5836 2540
rect 6836 1540 7046 2540
rect 5716 1487 7046 1540
rect 7134 1487 7196 2593
rect 5716 1420 7196 1487
rect 7330 2593 8810 2660
rect 7330 2540 8660 2593
rect 7330 1540 7450 2540
rect 8450 1540 8660 2540
rect 7330 1487 8660 1540
rect 8748 1487 8810 2593
rect 7330 1420 8810 1487
rect -8810 1233 -7330 1300
rect -8810 1180 -7480 1233
rect -8810 180 -8690 1180
rect -7690 180 -7480 1180
rect -8810 127 -7480 180
rect -7392 127 -7330 1233
rect -8810 60 -7330 127
rect -7196 1233 -5716 1300
rect -7196 1180 -5866 1233
rect -7196 180 -7076 1180
rect -6076 180 -5866 1180
rect -7196 127 -5866 180
rect -5778 127 -5716 1233
rect -7196 60 -5716 127
rect -5582 1233 -4102 1300
rect -5582 1180 -4252 1233
rect -5582 180 -5462 1180
rect -4462 180 -4252 1180
rect -5582 127 -4252 180
rect -4164 127 -4102 1233
rect -5582 60 -4102 127
rect -3968 1233 -2488 1300
rect -3968 1180 -2638 1233
rect -3968 180 -3848 1180
rect -2848 180 -2638 1180
rect -3968 127 -2638 180
rect -2550 127 -2488 1233
rect -3968 60 -2488 127
rect -2354 1233 -874 1300
rect -2354 1180 -1024 1233
rect -2354 180 -2234 1180
rect -1234 180 -1024 1180
rect -2354 127 -1024 180
rect -936 127 -874 1233
rect -2354 60 -874 127
rect -740 1233 740 1300
rect -740 1180 590 1233
rect -740 180 -620 1180
rect 380 180 590 1180
rect -740 127 590 180
rect 678 127 740 1233
rect -740 60 740 127
rect 874 1233 2354 1300
rect 874 1180 2204 1233
rect 874 180 994 1180
rect 1994 180 2204 1180
rect 874 127 2204 180
rect 2292 127 2354 1233
rect 874 60 2354 127
rect 2488 1233 3968 1300
rect 2488 1180 3818 1233
rect 2488 180 2608 1180
rect 3608 180 3818 1180
rect 2488 127 3818 180
rect 3906 127 3968 1233
rect 2488 60 3968 127
rect 4102 1233 5582 1300
rect 4102 1180 5432 1233
rect 4102 180 4222 1180
rect 5222 180 5432 1180
rect 4102 127 5432 180
rect 5520 127 5582 1233
rect 4102 60 5582 127
rect 5716 1233 7196 1300
rect 5716 1180 7046 1233
rect 5716 180 5836 1180
rect 6836 180 7046 1180
rect 5716 127 7046 180
rect 7134 127 7196 1233
rect 5716 60 7196 127
rect 7330 1233 8810 1300
rect 7330 1180 8660 1233
rect 7330 180 7450 1180
rect 8450 180 8660 1180
rect 7330 127 8660 180
rect 8748 127 8810 1233
rect 7330 60 8810 127
rect -8810 -127 -7330 -60
rect -8810 -180 -7480 -127
rect -8810 -1180 -8690 -180
rect -7690 -1180 -7480 -180
rect -8810 -1233 -7480 -1180
rect -7392 -1233 -7330 -127
rect -8810 -1300 -7330 -1233
rect -7196 -127 -5716 -60
rect -7196 -180 -5866 -127
rect -7196 -1180 -7076 -180
rect -6076 -1180 -5866 -180
rect -7196 -1233 -5866 -1180
rect -5778 -1233 -5716 -127
rect -7196 -1300 -5716 -1233
rect -5582 -127 -4102 -60
rect -5582 -180 -4252 -127
rect -5582 -1180 -5462 -180
rect -4462 -1180 -4252 -180
rect -5582 -1233 -4252 -1180
rect -4164 -1233 -4102 -127
rect -5582 -1300 -4102 -1233
rect -3968 -127 -2488 -60
rect -3968 -180 -2638 -127
rect -3968 -1180 -3848 -180
rect -2848 -1180 -2638 -180
rect -3968 -1233 -2638 -1180
rect -2550 -1233 -2488 -127
rect -3968 -1300 -2488 -1233
rect -2354 -127 -874 -60
rect -2354 -180 -1024 -127
rect -2354 -1180 -2234 -180
rect -1234 -1180 -1024 -180
rect -2354 -1233 -1024 -1180
rect -936 -1233 -874 -127
rect -2354 -1300 -874 -1233
rect -740 -127 740 -60
rect -740 -180 590 -127
rect -740 -1180 -620 -180
rect 380 -1180 590 -180
rect -740 -1233 590 -1180
rect 678 -1233 740 -127
rect -740 -1300 740 -1233
rect 874 -127 2354 -60
rect 874 -180 2204 -127
rect 874 -1180 994 -180
rect 1994 -1180 2204 -180
rect 874 -1233 2204 -1180
rect 2292 -1233 2354 -127
rect 874 -1300 2354 -1233
rect 2488 -127 3968 -60
rect 2488 -180 3818 -127
rect 2488 -1180 2608 -180
rect 3608 -1180 3818 -180
rect 2488 -1233 3818 -1180
rect 3906 -1233 3968 -127
rect 2488 -1300 3968 -1233
rect 4102 -127 5582 -60
rect 4102 -180 5432 -127
rect 4102 -1180 4222 -180
rect 5222 -1180 5432 -180
rect 4102 -1233 5432 -1180
rect 5520 -1233 5582 -127
rect 4102 -1300 5582 -1233
rect 5716 -127 7196 -60
rect 5716 -180 7046 -127
rect 5716 -1180 5836 -180
rect 6836 -1180 7046 -180
rect 5716 -1233 7046 -1180
rect 7134 -1233 7196 -127
rect 5716 -1300 7196 -1233
rect 7330 -127 8810 -60
rect 7330 -180 8660 -127
rect 7330 -1180 7450 -180
rect 8450 -1180 8660 -180
rect 7330 -1233 8660 -1180
rect 8748 -1233 8810 -127
rect 7330 -1300 8810 -1233
rect -8810 -1487 -7330 -1420
rect -8810 -1540 -7480 -1487
rect -8810 -2540 -8690 -1540
rect -7690 -2540 -7480 -1540
rect -8810 -2593 -7480 -2540
rect -7392 -2593 -7330 -1487
rect -8810 -2660 -7330 -2593
rect -7196 -1487 -5716 -1420
rect -7196 -1540 -5866 -1487
rect -7196 -2540 -7076 -1540
rect -6076 -2540 -5866 -1540
rect -7196 -2593 -5866 -2540
rect -5778 -2593 -5716 -1487
rect -7196 -2660 -5716 -2593
rect -5582 -1487 -4102 -1420
rect -5582 -1540 -4252 -1487
rect -5582 -2540 -5462 -1540
rect -4462 -2540 -4252 -1540
rect -5582 -2593 -4252 -2540
rect -4164 -2593 -4102 -1487
rect -5582 -2660 -4102 -2593
rect -3968 -1487 -2488 -1420
rect -3968 -1540 -2638 -1487
rect -3968 -2540 -3848 -1540
rect -2848 -2540 -2638 -1540
rect -3968 -2593 -2638 -2540
rect -2550 -2593 -2488 -1487
rect -3968 -2660 -2488 -2593
rect -2354 -1487 -874 -1420
rect -2354 -1540 -1024 -1487
rect -2354 -2540 -2234 -1540
rect -1234 -2540 -1024 -1540
rect -2354 -2593 -1024 -2540
rect -936 -2593 -874 -1487
rect -2354 -2660 -874 -2593
rect -740 -1487 740 -1420
rect -740 -1540 590 -1487
rect -740 -2540 -620 -1540
rect 380 -2540 590 -1540
rect -740 -2593 590 -2540
rect 678 -2593 740 -1487
rect -740 -2660 740 -2593
rect 874 -1487 2354 -1420
rect 874 -1540 2204 -1487
rect 874 -2540 994 -1540
rect 1994 -2540 2204 -1540
rect 874 -2593 2204 -2540
rect 2292 -2593 2354 -1487
rect 874 -2660 2354 -2593
rect 2488 -1487 3968 -1420
rect 2488 -1540 3818 -1487
rect 2488 -2540 2608 -1540
rect 3608 -2540 3818 -1540
rect 2488 -2593 3818 -2540
rect 3906 -2593 3968 -1487
rect 2488 -2660 3968 -2593
rect 4102 -1487 5582 -1420
rect 4102 -1540 5432 -1487
rect 4102 -2540 4222 -1540
rect 5222 -2540 5432 -1540
rect 4102 -2593 5432 -2540
rect 5520 -2593 5582 -1487
rect 4102 -2660 5582 -2593
rect 5716 -1487 7196 -1420
rect 5716 -1540 7046 -1487
rect 5716 -2540 5836 -1540
rect 6836 -2540 7046 -1540
rect 5716 -2593 7046 -2540
rect 7134 -2593 7196 -1487
rect 5716 -2660 7196 -2593
rect 7330 -1487 8810 -1420
rect 7330 -1540 8660 -1487
rect 7330 -2540 7450 -1540
rect 8450 -2540 8660 -1540
rect 7330 -2593 8660 -2540
rect 8748 -2593 8810 -1487
rect 7330 -2660 8810 -2593
rect -8810 -2847 -7330 -2780
rect -8810 -2900 -7480 -2847
rect -8810 -3900 -8690 -2900
rect -7690 -3900 -7480 -2900
rect -8810 -3953 -7480 -3900
rect -7392 -3953 -7330 -2847
rect -8810 -4020 -7330 -3953
rect -7196 -2847 -5716 -2780
rect -7196 -2900 -5866 -2847
rect -7196 -3900 -7076 -2900
rect -6076 -3900 -5866 -2900
rect -7196 -3953 -5866 -3900
rect -5778 -3953 -5716 -2847
rect -7196 -4020 -5716 -3953
rect -5582 -2847 -4102 -2780
rect -5582 -2900 -4252 -2847
rect -5582 -3900 -5462 -2900
rect -4462 -3900 -4252 -2900
rect -5582 -3953 -4252 -3900
rect -4164 -3953 -4102 -2847
rect -5582 -4020 -4102 -3953
rect -3968 -2847 -2488 -2780
rect -3968 -2900 -2638 -2847
rect -3968 -3900 -3848 -2900
rect -2848 -3900 -2638 -2900
rect -3968 -3953 -2638 -3900
rect -2550 -3953 -2488 -2847
rect -3968 -4020 -2488 -3953
rect -2354 -2847 -874 -2780
rect -2354 -2900 -1024 -2847
rect -2354 -3900 -2234 -2900
rect -1234 -3900 -1024 -2900
rect -2354 -3953 -1024 -3900
rect -936 -3953 -874 -2847
rect -2354 -4020 -874 -3953
rect -740 -2847 740 -2780
rect -740 -2900 590 -2847
rect -740 -3900 -620 -2900
rect 380 -3900 590 -2900
rect -740 -3953 590 -3900
rect 678 -3953 740 -2847
rect -740 -4020 740 -3953
rect 874 -2847 2354 -2780
rect 874 -2900 2204 -2847
rect 874 -3900 994 -2900
rect 1994 -3900 2204 -2900
rect 874 -3953 2204 -3900
rect 2292 -3953 2354 -2847
rect 874 -4020 2354 -3953
rect 2488 -2847 3968 -2780
rect 2488 -2900 3818 -2847
rect 2488 -3900 2608 -2900
rect 3608 -3900 3818 -2900
rect 2488 -3953 3818 -3900
rect 3906 -3953 3968 -2847
rect 2488 -4020 3968 -3953
rect 4102 -2847 5582 -2780
rect 4102 -2900 5432 -2847
rect 4102 -3900 4222 -2900
rect 5222 -3900 5432 -2900
rect 4102 -3953 5432 -3900
rect 5520 -3953 5582 -2847
rect 4102 -4020 5582 -3953
rect 5716 -2847 7196 -2780
rect 5716 -2900 7046 -2847
rect 5716 -3900 5836 -2900
rect 6836 -3900 7046 -2900
rect 5716 -3953 7046 -3900
rect 7134 -3953 7196 -2847
rect 5716 -4020 7196 -3953
rect 7330 -2847 8810 -2780
rect 7330 -2900 8660 -2847
rect 7330 -3900 7450 -2900
rect 8450 -3900 8660 -2900
rect 7330 -3953 8660 -3900
rect 8748 -3953 8810 -2847
rect 7330 -4020 8810 -3953
rect -8810 -4207 -7330 -4140
rect -8810 -4260 -7480 -4207
rect -8810 -5260 -8690 -4260
rect -7690 -5260 -7480 -4260
rect -8810 -5313 -7480 -5260
rect -7392 -5313 -7330 -4207
rect -8810 -5380 -7330 -5313
rect -7196 -4207 -5716 -4140
rect -7196 -4260 -5866 -4207
rect -7196 -5260 -7076 -4260
rect -6076 -5260 -5866 -4260
rect -7196 -5313 -5866 -5260
rect -5778 -5313 -5716 -4207
rect -7196 -5380 -5716 -5313
rect -5582 -4207 -4102 -4140
rect -5582 -4260 -4252 -4207
rect -5582 -5260 -5462 -4260
rect -4462 -5260 -4252 -4260
rect -5582 -5313 -4252 -5260
rect -4164 -5313 -4102 -4207
rect -5582 -5380 -4102 -5313
rect -3968 -4207 -2488 -4140
rect -3968 -4260 -2638 -4207
rect -3968 -5260 -3848 -4260
rect -2848 -5260 -2638 -4260
rect -3968 -5313 -2638 -5260
rect -2550 -5313 -2488 -4207
rect -3968 -5380 -2488 -5313
rect -2354 -4207 -874 -4140
rect -2354 -4260 -1024 -4207
rect -2354 -5260 -2234 -4260
rect -1234 -5260 -1024 -4260
rect -2354 -5313 -1024 -5260
rect -936 -5313 -874 -4207
rect -2354 -5380 -874 -5313
rect -740 -4207 740 -4140
rect -740 -4260 590 -4207
rect -740 -5260 -620 -4260
rect 380 -5260 590 -4260
rect -740 -5313 590 -5260
rect 678 -5313 740 -4207
rect -740 -5380 740 -5313
rect 874 -4207 2354 -4140
rect 874 -4260 2204 -4207
rect 874 -5260 994 -4260
rect 1994 -5260 2204 -4260
rect 874 -5313 2204 -5260
rect 2292 -5313 2354 -4207
rect 874 -5380 2354 -5313
rect 2488 -4207 3968 -4140
rect 2488 -4260 3818 -4207
rect 2488 -5260 2608 -4260
rect 3608 -5260 3818 -4260
rect 2488 -5313 3818 -5260
rect 3906 -5313 3968 -4207
rect 2488 -5380 3968 -5313
rect 4102 -4207 5582 -4140
rect 4102 -4260 5432 -4207
rect 4102 -5260 4222 -4260
rect 5222 -5260 5432 -4260
rect 4102 -5313 5432 -5260
rect 5520 -5313 5582 -4207
rect 4102 -5380 5582 -5313
rect 5716 -4207 7196 -4140
rect 5716 -4260 7046 -4207
rect 5716 -5260 5836 -4260
rect 6836 -5260 7046 -4260
rect 5716 -5313 7046 -5260
rect 7134 -5313 7196 -4207
rect 5716 -5380 7196 -5313
rect 7330 -4207 8810 -4140
rect 7330 -4260 8660 -4207
rect 7330 -5260 7450 -4260
rect 8450 -5260 8660 -4260
rect 7330 -5313 8660 -5260
rect 8748 -5313 8810 -4207
rect 7330 -5380 8810 -5313
rect -8810 -5567 -7330 -5500
rect -8810 -5620 -7480 -5567
rect -8810 -6620 -8690 -5620
rect -7690 -6620 -7480 -5620
rect -8810 -6673 -7480 -6620
rect -7392 -6673 -7330 -5567
rect -8810 -6740 -7330 -6673
rect -7196 -5567 -5716 -5500
rect -7196 -5620 -5866 -5567
rect -7196 -6620 -7076 -5620
rect -6076 -6620 -5866 -5620
rect -7196 -6673 -5866 -6620
rect -5778 -6673 -5716 -5567
rect -7196 -6740 -5716 -6673
rect -5582 -5567 -4102 -5500
rect -5582 -5620 -4252 -5567
rect -5582 -6620 -5462 -5620
rect -4462 -6620 -4252 -5620
rect -5582 -6673 -4252 -6620
rect -4164 -6673 -4102 -5567
rect -5582 -6740 -4102 -6673
rect -3968 -5567 -2488 -5500
rect -3968 -5620 -2638 -5567
rect -3968 -6620 -3848 -5620
rect -2848 -6620 -2638 -5620
rect -3968 -6673 -2638 -6620
rect -2550 -6673 -2488 -5567
rect -3968 -6740 -2488 -6673
rect -2354 -5567 -874 -5500
rect -2354 -5620 -1024 -5567
rect -2354 -6620 -2234 -5620
rect -1234 -6620 -1024 -5620
rect -2354 -6673 -1024 -6620
rect -936 -6673 -874 -5567
rect -2354 -6740 -874 -6673
rect -740 -5567 740 -5500
rect -740 -5620 590 -5567
rect -740 -6620 -620 -5620
rect 380 -6620 590 -5620
rect -740 -6673 590 -6620
rect 678 -6673 740 -5567
rect -740 -6740 740 -6673
rect 874 -5567 2354 -5500
rect 874 -5620 2204 -5567
rect 874 -6620 994 -5620
rect 1994 -6620 2204 -5620
rect 874 -6673 2204 -6620
rect 2292 -6673 2354 -5567
rect 874 -6740 2354 -6673
rect 2488 -5567 3968 -5500
rect 2488 -5620 3818 -5567
rect 2488 -6620 2608 -5620
rect 3608 -6620 3818 -5620
rect 2488 -6673 3818 -6620
rect 3906 -6673 3968 -5567
rect 2488 -6740 3968 -6673
rect 4102 -5567 5582 -5500
rect 4102 -5620 5432 -5567
rect 4102 -6620 4222 -5620
rect 5222 -6620 5432 -5620
rect 4102 -6673 5432 -6620
rect 5520 -6673 5582 -5567
rect 4102 -6740 5582 -6673
rect 5716 -5567 7196 -5500
rect 5716 -5620 7046 -5567
rect 5716 -6620 5836 -5620
rect 6836 -6620 7046 -5620
rect 5716 -6673 7046 -6620
rect 7134 -6673 7196 -5567
rect 5716 -6740 7196 -6673
rect 7330 -5567 8810 -5500
rect 7330 -5620 8660 -5567
rect 7330 -6620 7450 -5620
rect 8450 -6620 8660 -5620
rect 7330 -6673 8660 -6620
rect 8748 -6673 8810 -5567
rect 7330 -6740 8810 -6673
rect -8810 -6927 -7330 -6860
rect -8810 -6980 -7480 -6927
rect -8810 -7980 -8690 -6980
rect -7690 -7980 -7480 -6980
rect -8810 -8033 -7480 -7980
rect -7392 -8033 -7330 -6927
rect -8810 -8100 -7330 -8033
rect -7196 -6927 -5716 -6860
rect -7196 -6980 -5866 -6927
rect -7196 -7980 -7076 -6980
rect -6076 -7980 -5866 -6980
rect -7196 -8033 -5866 -7980
rect -5778 -8033 -5716 -6927
rect -7196 -8100 -5716 -8033
rect -5582 -6927 -4102 -6860
rect -5582 -6980 -4252 -6927
rect -5582 -7980 -5462 -6980
rect -4462 -7980 -4252 -6980
rect -5582 -8033 -4252 -7980
rect -4164 -8033 -4102 -6927
rect -5582 -8100 -4102 -8033
rect -3968 -6927 -2488 -6860
rect -3968 -6980 -2638 -6927
rect -3968 -7980 -3848 -6980
rect -2848 -7980 -2638 -6980
rect -3968 -8033 -2638 -7980
rect -2550 -8033 -2488 -6927
rect -3968 -8100 -2488 -8033
rect -2354 -6927 -874 -6860
rect -2354 -6980 -1024 -6927
rect -2354 -7980 -2234 -6980
rect -1234 -7980 -1024 -6980
rect -2354 -8033 -1024 -7980
rect -936 -8033 -874 -6927
rect -2354 -8100 -874 -8033
rect -740 -6927 740 -6860
rect -740 -6980 590 -6927
rect -740 -7980 -620 -6980
rect 380 -7980 590 -6980
rect -740 -8033 590 -7980
rect 678 -8033 740 -6927
rect -740 -8100 740 -8033
rect 874 -6927 2354 -6860
rect 874 -6980 2204 -6927
rect 874 -7980 994 -6980
rect 1994 -7980 2204 -6980
rect 874 -8033 2204 -7980
rect 2292 -8033 2354 -6927
rect 874 -8100 2354 -8033
rect 2488 -6927 3968 -6860
rect 2488 -6980 3818 -6927
rect 2488 -7980 2608 -6980
rect 3608 -7980 3818 -6980
rect 2488 -8033 3818 -7980
rect 3906 -8033 3968 -6927
rect 2488 -8100 3968 -8033
rect 4102 -6927 5582 -6860
rect 4102 -6980 5432 -6927
rect 4102 -7980 4222 -6980
rect 5222 -7980 5432 -6980
rect 4102 -8033 5432 -7980
rect 5520 -8033 5582 -6927
rect 4102 -8100 5582 -8033
rect 5716 -6927 7196 -6860
rect 5716 -6980 7046 -6927
rect 5716 -7980 5836 -6980
rect 6836 -7980 7046 -6980
rect 5716 -8033 7046 -7980
rect 7134 -8033 7196 -6927
rect 5716 -8100 7196 -8033
rect 7330 -6927 8810 -6860
rect 7330 -6980 8660 -6927
rect 7330 -7980 7450 -6980
rect 8450 -7980 8660 -6980
rect 7330 -8033 8660 -7980
rect 8748 -8033 8810 -6927
rect 7330 -8100 8810 -8033
<< via4 >>
rect -7480 6927 -7392 8033
rect -5866 6927 -5778 8033
rect -4252 6927 -4164 8033
rect -2638 6927 -2550 8033
rect -1024 6927 -936 8033
rect 590 6927 678 8033
rect 2204 6927 2292 8033
rect 3818 6927 3906 8033
rect 5432 6927 5520 8033
rect 7046 6927 7134 8033
rect 8660 6927 8748 8033
rect -7480 5567 -7392 6673
rect -5866 5567 -5778 6673
rect -4252 5567 -4164 6673
rect -2638 5567 -2550 6673
rect -1024 5567 -936 6673
rect 590 5567 678 6673
rect 2204 5567 2292 6673
rect 3818 5567 3906 6673
rect 5432 5567 5520 6673
rect 7046 5567 7134 6673
rect 8660 5567 8748 6673
rect -7480 4207 -7392 5313
rect -5866 4207 -5778 5313
rect -4252 4207 -4164 5313
rect -2638 4207 -2550 5313
rect -1024 4207 -936 5313
rect 590 4207 678 5313
rect 2204 4207 2292 5313
rect 3818 4207 3906 5313
rect 5432 4207 5520 5313
rect 7046 4207 7134 5313
rect 8660 4207 8748 5313
rect -7480 2847 -7392 3953
rect -5866 2847 -5778 3953
rect -4252 2847 -4164 3953
rect -2638 2847 -2550 3953
rect -1024 2847 -936 3953
rect 590 2847 678 3953
rect 2204 2847 2292 3953
rect 3818 2847 3906 3953
rect 5432 2847 5520 3953
rect 7046 2847 7134 3953
rect 8660 2847 8748 3953
rect -7480 1487 -7392 2593
rect -5866 1487 -5778 2593
rect -4252 1487 -4164 2593
rect -2638 1487 -2550 2593
rect -1024 1487 -936 2593
rect 590 1487 678 2593
rect 2204 1487 2292 2593
rect 3818 1487 3906 2593
rect 5432 1487 5520 2593
rect 7046 1487 7134 2593
rect 8660 1487 8748 2593
rect -7480 127 -7392 1233
rect -5866 127 -5778 1233
rect -4252 127 -4164 1233
rect -2638 127 -2550 1233
rect -1024 127 -936 1233
rect 590 127 678 1233
rect 2204 127 2292 1233
rect 3818 127 3906 1233
rect 5432 127 5520 1233
rect 7046 127 7134 1233
rect 8660 127 8748 1233
rect -7480 -1233 -7392 -127
rect -5866 -1233 -5778 -127
rect -4252 -1233 -4164 -127
rect -2638 -1233 -2550 -127
rect -1024 -1233 -936 -127
rect 590 -1233 678 -127
rect 2204 -1233 2292 -127
rect 3818 -1233 3906 -127
rect 5432 -1233 5520 -127
rect 7046 -1233 7134 -127
rect 8660 -1233 8748 -127
rect -7480 -2593 -7392 -1487
rect -5866 -2593 -5778 -1487
rect -4252 -2593 -4164 -1487
rect -2638 -2593 -2550 -1487
rect -1024 -2593 -936 -1487
rect 590 -2593 678 -1487
rect 2204 -2593 2292 -1487
rect 3818 -2593 3906 -1487
rect 5432 -2593 5520 -1487
rect 7046 -2593 7134 -1487
rect 8660 -2593 8748 -1487
rect -7480 -3953 -7392 -2847
rect -5866 -3953 -5778 -2847
rect -4252 -3953 -4164 -2847
rect -2638 -3953 -2550 -2847
rect -1024 -3953 -936 -2847
rect 590 -3953 678 -2847
rect 2204 -3953 2292 -2847
rect 3818 -3953 3906 -2847
rect 5432 -3953 5520 -2847
rect 7046 -3953 7134 -2847
rect 8660 -3953 8748 -2847
rect -7480 -5313 -7392 -4207
rect -5866 -5313 -5778 -4207
rect -4252 -5313 -4164 -4207
rect -2638 -5313 -2550 -4207
rect -1024 -5313 -936 -4207
rect 590 -5313 678 -4207
rect 2204 -5313 2292 -4207
rect 3818 -5313 3906 -4207
rect 5432 -5313 5520 -4207
rect 7046 -5313 7134 -4207
rect 8660 -5313 8748 -4207
rect -7480 -6673 -7392 -5567
rect -5866 -6673 -5778 -5567
rect -4252 -6673 -4164 -5567
rect -2638 -6673 -2550 -5567
rect -1024 -6673 -936 -5567
rect 590 -6673 678 -5567
rect 2204 -6673 2292 -5567
rect 3818 -6673 3906 -5567
rect 5432 -6673 5520 -5567
rect 7046 -6673 7134 -5567
rect 8660 -6673 8748 -5567
rect -7480 -8033 -7392 -6927
rect -5866 -8033 -5778 -6927
rect -4252 -8033 -4164 -6927
rect -2638 -8033 -2550 -6927
rect -1024 -8033 -936 -6927
rect 590 -8033 678 -6927
rect 2204 -8033 2292 -6927
rect 3818 -8033 3906 -6927
rect 5432 -8033 5520 -6927
rect 7046 -8033 7134 -6927
rect 8660 -8033 8748 -6927
<< metal5 >>
rect -8296 7900 -8084 8160
rect -7542 8033 -7330 8160
rect -8296 6540 -8084 7060
rect -7542 6927 -7480 8033
rect -7392 6927 -7330 8033
rect -6682 7900 -6470 8160
rect -5928 8033 -5716 8160
rect -7542 6673 -7330 6927
rect -8296 5180 -8084 5700
rect -7542 5567 -7480 6673
rect -7392 5567 -7330 6673
rect -6682 6540 -6470 7060
rect -5928 6927 -5866 8033
rect -5778 6927 -5716 8033
rect -5068 7900 -4856 8160
rect -4314 8033 -4102 8160
rect -5928 6673 -5716 6927
rect -7542 5313 -7330 5567
rect -8296 3820 -8084 4340
rect -7542 4207 -7480 5313
rect -7392 4207 -7330 5313
rect -6682 5180 -6470 5700
rect -5928 5567 -5866 6673
rect -5778 5567 -5716 6673
rect -5068 6540 -4856 7060
rect -4314 6927 -4252 8033
rect -4164 6927 -4102 8033
rect -3454 7900 -3242 8160
rect -2700 8033 -2488 8160
rect -4314 6673 -4102 6927
rect -5928 5313 -5716 5567
rect -7542 3953 -7330 4207
rect -8296 2460 -8084 2980
rect -7542 2847 -7480 3953
rect -7392 2847 -7330 3953
rect -6682 3820 -6470 4340
rect -5928 4207 -5866 5313
rect -5778 4207 -5716 5313
rect -5068 5180 -4856 5700
rect -4314 5567 -4252 6673
rect -4164 5567 -4102 6673
rect -3454 6540 -3242 7060
rect -2700 6927 -2638 8033
rect -2550 6927 -2488 8033
rect -1840 7900 -1628 8160
rect -1086 8033 -874 8160
rect -2700 6673 -2488 6927
rect -4314 5313 -4102 5567
rect -5928 3953 -5716 4207
rect -7542 2593 -7330 2847
rect -8296 1100 -8084 1620
rect -7542 1487 -7480 2593
rect -7392 1487 -7330 2593
rect -6682 2460 -6470 2980
rect -5928 2847 -5866 3953
rect -5778 2847 -5716 3953
rect -5068 3820 -4856 4340
rect -4314 4207 -4252 5313
rect -4164 4207 -4102 5313
rect -3454 5180 -3242 5700
rect -2700 5567 -2638 6673
rect -2550 5567 -2488 6673
rect -1840 6540 -1628 7060
rect -1086 6927 -1024 8033
rect -936 6927 -874 8033
rect -226 7900 -14 8160
rect 528 8033 740 8160
rect -1086 6673 -874 6927
rect -2700 5313 -2488 5567
rect -4314 3953 -4102 4207
rect -5928 2593 -5716 2847
rect -7542 1233 -7330 1487
rect -8296 -260 -8084 260
rect -7542 127 -7480 1233
rect -7392 127 -7330 1233
rect -6682 1100 -6470 1620
rect -5928 1487 -5866 2593
rect -5778 1487 -5716 2593
rect -5068 2460 -4856 2980
rect -4314 2847 -4252 3953
rect -4164 2847 -4102 3953
rect -3454 3820 -3242 4340
rect -2700 4207 -2638 5313
rect -2550 4207 -2488 5313
rect -1840 5180 -1628 5700
rect -1086 5567 -1024 6673
rect -936 5567 -874 6673
rect -226 6540 -14 7060
rect 528 6927 590 8033
rect 678 6927 740 8033
rect 1388 7900 1600 8160
rect 2142 8033 2354 8160
rect 528 6673 740 6927
rect -1086 5313 -874 5567
rect -2700 3953 -2488 4207
rect -4314 2593 -4102 2847
rect -5928 1233 -5716 1487
rect -7542 -127 -7330 127
rect -8296 -1620 -8084 -1100
rect -7542 -1233 -7480 -127
rect -7392 -1233 -7330 -127
rect -6682 -260 -6470 260
rect -5928 127 -5866 1233
rect -5778 127 -5716 1233
rect -5068 1100 -4856 1620
rect -4314 1487 -4252 2593
rect -4164 1487 -4102 2593
rect -3454 2460 -3242 2980
rect -2700 2847 -2638 3953
rect -2550 2847 -2488 3953
rect -1840 3820 -1628 4340
rect -1086 4207 -1024 5313
rect -936 4207 -874 5313
rect -226 5180 -14 5700
rect 528 5567 590 6673
rect 678 5567 740 6673
rect 1388 6540 1600 7060
rect 2142 6927 2204 8033
rect 2292 6927 2354 8033
rect 3002 7900 3214 8160
rect 3756 8033 3968 8160
rect 2142 6673 2354 6927
rect 528 5313 740 5567
rect -1086 3953 -874 4207
rect -2700 2593 -2488 2847
rect -4314 1233 -4102 1487
rect -5928 -127 -5716 127
rect -7542 -1487 -7330 -1233
rect -8296 -2980 -8084 -2460
rect -7542 -2593 -7480 -1487
rect -7392 -2593 -7330 -1487
rect -6682 -1620 -6470 -1100
rect -5928 -1233 -5866 -127
rect -5778 -1233 -5716 -127
rect -5068 -260 -4856 260
rect -4314 127 -4252 1233
rect -4164 127 -4102 1233
rect -3454 1100 -3242 1620
rect -2700 1487 -2638 2593
rect -2550 1487 -2488 2593
rect -1840 2460 -1628 2980
rect -1086 2847 -1024 3953
rect -936 2847 -874 3953
rect -226 3820 -14 4340
rect 528 4207 590 5313
rect 678 4207 740 5313
rect 1388 5180 1600 5700
rect 2142 5567 2204 6673
rect 2292 5567 2354 6673
rect 3002 6540 3214 7060
rect 3756 6927 3818 8033
rect 3906 6927 3968 8033
rect 4616 7900 4828 8160
rect 5370 8033 5582 8160
rect 3756 6673 3968 6927
rect 2142 5313 2354 5567
rect 528 3953 740 4207
rect -1086 2593 -874 2847
rect -2700 1233 -2488 1487
rect -4314 -127 -4102 127
rect -5928 -1487 -5716 -1233
rect -7542 -2847 -7330 -2593
rect -8296 -4340 -8084 -3820
rect -7542 -3953 -7480 -2847
rect -7392 -3953 -7330 -2847
rect -6682 -2980 -6470 -2460
rect -5928 -2593 -5866 -1487
rect -5778 -2593 -5716 -1487
rect -5068 -1620 -4856 -1100
rect -4314 -1233 -4252 -127
rect -4164 -1233 -4102 -127
rect -3454 -260 -3242 260
rect -2700 127 -2638 1233
rect -2550 127 -2488 1233
rect -1840 1100 -1628 1620
rect -1086 1487 -1024 2593
rect -936 1487 -874 2593
rect -226 2460 -14 2980
rect 528 2847 590 3953
rect 678 2847 740 3953
rect 1388 3820 1600 4340
rect 2142 4207 2204 5313
rect 2292 4207 2354 5313
rect 3002 5180 3214 5700
rect 3756 5567 3818 6673
rect 3906 5567 3968 6673
rect 4616 6540 4828 7060
rect 5370 6927 5432 8033
rect 5520 6927 5582 8033
rect 6230 7900 6442 8160
rect 6984 8033 7196 8160
rect 5370 6673 5582 6927
rect 3756 5313 3968 5567
rect 2142 3953 2354 4207
rect 528 2593 740 2847
rect -1086 1233 -874 1487
rect -2700 -127 -2488 127
rect -4314 -1487 -4102 -1233
rect -5928 -2847 -5716 -2593
rect -7542 -4207 -7330 -3953
rect -8296 -5700 -8084 -5180
rect -7542 -5313 -7480 -4207
rect -7392 -5313 -7330 -4207
rect -6682 -4340 -6470 -3820
rect -5928 -3953 -5866 -2847
rect -5778 -3953 -5716 -2847
rect -5068 -2980 -4856 -2460
rect -4314 -2593 -4252 -1487
rect -4164 -2593 -4102 -1487
rect -3454 -1620 -3242 -1100
rect -2700 -1233 -2638 -127
rect -2550 -1233 -2488 -127
rect -1840 -260 -1628 260
rect -1086 127 -1024 1233
rect -936 127 -874 1233
rect -226 1100 -14 1620
rect 528 1487 590 2593
rect 678 1487 740 2593
rect 1388 2460 1600 2980
rect 2142 2847 2204 3953
rect 2292 2847 2354 3953
rect 3002 3820 3214 4340
rect 3756 4207 3818 5313
rect 3906 4207 3968 5313
rect 4616 5180 4828 5700
rect 5370 5567 5432 6673
rect 5520 5567 5582 6673
rect 6230 6540 6442 7060
rect 6984 6927 7046 8033
rect 7134 6927 7196 8033
rect 7844 7900 8056 8160
rect 8598 8033 8810 8160
rect 6984 6673 7196 6927
rect 5370 5313 5582 5567
rect 3756 3953 3968 4207
rect 2142 2593 2354 2847
rect 528 1233 740 1487
rect -1086 -127 -874 127
rect -2700 -1487 -2488 -1233
rect -4314 -2847 -4102 -2593
rect -5928 -4207 -5716 -3953
rect -7542 -5567 -7330 -5313
rect -8296 -7060 -8084 -6540
rect -7542 -6673 -7480 -5567
rect -7392 -6673 -7330 -5567
rect -6682 -5700 -6470 -5180
rect -5928 -5313 -5866 -4207
rect -5778 -5313 -5716 -4207
rect -5068 -4340 -4856 -3820
rect -4314 -3953 -4252 -2847
rect -4164 -3953 -4102 -2847
rect -3454 -2980 -3242 -2460
rect -2700 -2593 -2638 -1487
rect -2550 -2593 -2488 -1487
rect -1840 -1620 -1628 -1100
rect -1086 -1233 -1024 -127
rect -936 -1233 -874 -127
rect -226 -260 -14 260
rect 528 127 590 1233
rect 678 127 740 1233
rect 1388 1100 1600 1620
rect 2142 1487 2204 2593
rect 2292 1487 2354 2593
rect 3002 2460 3214 2980
rect 3756 2847 3818 3953
rect 3906 2847 3968 3953
rect 4616 3820 4828 4340
rect 5370 4207 5432 5313
rect 5520 4207 5582 5313
rect 6230 5180 6442 5700
rect 6984 5567 7046 6673
rect 7134 5567 7196 6673
rect 7844 6540 8056 7060
rect 8598 6927 8660 8033
rect 8748 6927 8810 8033
rect 8598 6673 8810 6927
rect 6984 5313 7196 5567
rect 5370 3953 5582 4207
rect 3756 2593 3968 2847
rect 2142 1233 2354 1487
rect 528 -127 740 127
rect -1086 -1487 -874 -1233
rect -2700 -2847 -2488 -2593
rect -4314 -4207 -4102 -3953
rect -5928 -5567 -5716 -5313
rect -7542 -6927 -7330 -6673
rect -8296 -8160 -8084 -7900
rect -7542 -8033 -7480 -6927
rect -7392 -8033 -7330 -6927
rect -6682 -7060 -6470 -6540
rect -5928 -6673 -5866 -5567
rect -5778 -6673 -5716 -5567
rect -5068 -5700 -4856 -5180
rect -4314 -5313 -4252 -4207
rect -4164 -5313 -4102 -4207
rect -3454 -4340 -3242 -3820
rect -2700 -3953 -2638 -2847
rect -2550 -3953 -2488 -2847
rect -1840 -2980 -1628 -2460
rect -1086 -2593 -1024 -1487
rect -936 -2593 -874 -1487
rect -226 -1620 -14 -1100
rect 528 -1233 590 -127
rect 678 -1233 740 -127
rect 1388 -260 1600 260
rect 2142 127 2204 1233
rect 2292 127 2354 1233
rect 3002 1100 3214 1620
rect 3756 1487 3818 2593
rect 3906 1487 3968 2593
rect 4616 2460 4828 2980
rect 5370 2847 5432 3953
rect 5520 2847 5582 3953
rect 6230 3820 6442 4340
rect 6984 4207 7046 5313
rect 7134 4207 7196 5313
rect 7844 5180 8056 5700
rect 8598 5567 8660 6673
rect 8748 5567 8810 6673
rect 8598 5313 8810 5567
rect 6984 3953 7196 4207
rect 5370 2593 5582 2847
rect 3756 1233 3968 1487
rect 2142 -127 2354 127
rect 528 -1487 740 -1233
rect -1086 -2847 -874 -2593
rect -2700 -4207 -2488 -3953
rect -4314 -5567 -4102 -5313
rect -5928 -6927 -5716 -6673
rect -7542 -8160 -7330 -8033
rect -6682 -8160 -6470 -7900
rect -5928 -8033 -5866 -6927
rect -5778 -8033 -5716 -6927
rect -5068 -7060 -4856 -6540
rect -4314 -6673 -4252 -5567
rect -4164 -6673 -4102 -5567
rect -3454 -5700 -3242 -5180
rect -2700 -5313 -2638 -4207
rect -2550 -5313 -2488 -4207
rect -1840 -4340 -1628 -3820
rect -1086 -3953 -1024 -2847
rect -936 -3953 -874 -2847
rect -226 -2980 -14 -2460
rect 528 -2593 590 -1487
rect 678 -2593 740 -1487
rect 1388 -1620 1600 -1100
rect 2142 -1233 2204 -127
rect 2292 -1233 2354 -127
rect 3002 -260 3214 260
rect 3756 127 3818 1233
rect 3906 127 3968 1233
rect 4616 1100 4828 1620
rect 5370 1487 5432 2593
rect 5520 1487 5582 2593
rect 6230 2460 6442 2980
rect 6984 2847 7046 3953
rect 7134 2847 7196 3953
rect 7844 3820 8056 4340
rect 8598 4207 8660 5313
rect 8748 4207 8810 5313
rect 8598 3953 8810 4207
rect 6984 2593 7196 2847
rect 5370 1233 5582 1487
rect 3756 -127 3968 127
rect 2142 -1487 2354 -1233
rect 528 -2847 740 -2593
rect -1086 -4207 -874 -3953
rect -2700 -5567 -2488 -5313
rect -4314 -6927 -4102 -6673
rect -5928 -8160 -5716 -8033
rect -5068 -8160 -4856 -7900
rect -4314 -8033 -4252 -6927
rect -4164 -8033 -4102 -6927
rect -3454 -7060 -3242 -6540
rect -2700 -6673 -2638 -5567
rect -2550 -6673 -2488 -5567
rect -1840 -5700 -1628 -5180
rect -1086 -5313 -1024 -4207
rect -936 -5313 -874 -4207
rect -226 -4340 -14 -3820
rect 528 -3953 590 -2847
rect 678 -3953 740 -2847
rect 1388 -2980 1600 -2460
rect 2142 -2593 2204 -1487
rect 2292 -2593 2354 -1487
rect 3002 -1620 3214 -1100
rect 3756 -1233 3818 -127
rect 3906 -1233 3968 -127
rect 4616 -260 4828 260
rect 5370 127 5432 1233
rect 5520 127 5582 1233
rect 6230 1100 6442 1620
rect 6984 1487 7046 2593
rect 7134 1487 7196 2593
rect 7844 2460 8056 2980
rect 8598 2847 8660 3953
rect 8748 2847 8810 3953
rect 8598 2593 8810 2847
rect 6984 1233 7196 1487
rect 5370 -127 5582 127
rect 3756 -1487 3968 -1233
rect 2142 -2847 2354 -2593
rect 528 -4207 740 -3953
rect -1086 -5567 -874 -5313
rect -2700 -6927 -2488 -6673
rect -4314 -8160 -4102 -8033
rect -3454 -8160 -3242 -7900
rect -2700 -8033 -2638 -6927
rect -2550 -8033 -2488 -6927
rect -1840 -7060 -1628 -6540
rect -1086 -6673 -1024 -5567
rect -936 -6673 -874 -5567
rect -226 -5700 -14 -5180
rect 528 -5313 590 -4207
rect 678 -5313 740 -4207
rect 1388 -4340 1600 -3820
rect 2142 -3953 2204 -2847
rect 2292 -3953 2354 -2847
rect 3002 -2980 3214 -2460
rect 3756 -2593 3818 -1487
rect 3906 -2593 3968 -1487
rect 4616 -1620 4828 -1100
rect 5370 -1233 5432 -127
rect 5520 -1233 5582 -127
rect 6230 -260 6442 260
rect 6984 127 7046 1233
rect 7134 127 7196 1233
rect 7844 1100 8056 1620
rect 8598 1487 8660 2593
rect 8748 1487 8810 2593
rect 8598 1233 8810 1487
rect 6984 -127 7196 127
rect 5370 -1487 5582 -1233
rect 3756 -2847 3968 -2593
rect 2142 -4207 2354 -3953
rect 528 -5567 740 -5313
rect -1086 -6927 -874 -6673
rect -2700 -8160 -2488 -8033
rect -1840 -8160 -1628 -7900
rect -1086 -8033 -1024 -6927
rect -936 -8033 -874 -6927
rect -226 -7060 -14 -6540
rect 528 -6673 590 -5567
rect 678 -6673 740 -5567
rect 1388 -5700 1600 -5180
rect 2142 -5313 2204 -4207
rect 2292 -5313 2354 -4207
rect 3002 -4340 3214 -3820
rect 3756 -3953 3818 -2847
rect 3906 -3953 3968 -2847
rect 4616 -2980 4828 -2460
rect 5370 -2593 5432 -1487
rect 5520 -2593 5582 -1487
rect 6230 -1620 6442 -1100
rect 6984 -1233 7046 -127
rect 7134 -1233 7196 -127
rect 7844 -260 8056 260
rect 8598 127 8660 1233
rect 8748 127 8810 1233
rect 8598 -127 8810 127
rect 6984 -1487 7196 -1233
rect 5370 -2847 5582 -2593
rect 3756 -4207 3968 -3953
rect 2142 -5567 2354 -5313
rect 528 -6927 740 -6673
rect -1086 -8160 -874 -8033
rect -226 -8160 -14 -7900
rect 528 -8033 590 -6927
rect 678 -8033 740 -6927
rect 1388 -7060 1600 -6540
rect 2142 -6673 2204 -5567
rect 2292 -6673 2354 -5567
rect 3002 -5700 3214 -5180
rect 3756 -5313 3818 -4207
rect 3906 -5313 3968 -4207
rect 4616 -4340 4828 -3820
rect 5370 -3953 5432 -2847
rect 5520 -3953 5582 -2847
rect 6230 -2980 6442 -2460
rect 6984 -2593 7046 -1487
rect 7134 -2593 7196 -1487
rect 7844 -1620 8056 -1100
rect 8598 -1233 8660 -127
rect 8748 -1233 8810 -127
rect 8598 -1487 8810 -1233
rect 6984 -2847 7196 -2593
rect 5370 -4207 5582 -3953
rect 3756 -5567 3968 -5313
rect 2142 -6927 2354 -6673
rect 528 -8160 740 -8033
rect 1388 -8160 1600 -7900
rect 2142 -8033 2204 -6927
rect 2292 -8033 2354 -6927
rect 3002 -7060 3214 -6540
rect 3756 -6673 3818 -5567
rect 3906 -6673 3968 -5567
rect 4616 -5700 4828 -5180
rect 5370 -5313 5432 -4207
rect 5520 -5313 5582 -4207
rect 6230 -4340 6442 -3820
rect 6984 -3953 7046 -2847
rect 7134 -3953 7196 -2847
rect 7844 -2980 8056 -2460
rect 8598 -2593 8660 -1487
rect 8748 -2593 8810 -1487
rect 8598 -2847 8810 -2593
rect 6984 -4207 7196 -3953
rect 5370 -5567 5582 -5313
rect 3756 -6927 3968 -6673
rect 2142 -8160 2354 -8033
rect 3002 -8160 3214 -7900
rect 3756 -8033 3818 -6927
rect 3906 -8033 3968 -6927
rect 4616 -7060 4828 -6540
rect 5370 -6673 5432 -5567
rect 5520 -6673 5582 -5567
rect 6230 -5700 6442 -5180
rect 6984 -5313 7046 -4207
rect 7134 -5313 7196 -4207
rect 7844 -4340 8056 -3820
rect 8598 -3953 8660 -2847
rect 8748 -3953 8810 -2847
rect 8598 -4207 8810 -3953
rect 6984 -5567 7196 -5313
rect 5370 -6927 5582 -6673
rect 3756 -8160 3968 -8033
rect 4616 -8160 4828 -7900
rect 5370 -8033 5432 -6927
rect 5520 -8033 5582 -6927
rect 6230 -7060 6442 -6540
rect 6984 -6673 7046 -5567
rect 7134 -6673 7196 -5567
rect 7844 -5700 8056 -5180
rect 8598 -5313 8660 -4207
rect 8748 -5313 8810 -4207
rect 8598 -5567 8810 -5313
rect 6984 -6927 7196 -6673
rect 5370 -8160 5582 -8033
rect 6230 -8160 6442 -7900
rect 6984 -8033 7046 -6927
rect 7134 -8033 7196 -6927
rect 7844 -7060 8056 -6540
rect 8598 -6673 8660 -5567
rect 8748 -6673 8810 -5567
rect 8598 -6927 8810 -6673
rect 6984 -8160 7196 -8033
rect 7844 -8160 8056 -7900
rect 8598 -8033 8660 -6927
rect 8748 -8033 8810 -6927
rect 8598 -8160 8810 -8033
<< properties >>
string FIXED_BBOX 7330 6860 8570 8100
string gencell cap_mim_2p0fF
string library gf180mcu
string parameters w 5.00 l 5.00 val 1.025k carea 25.00 cperi 20.00 class capacitor nx 11 ny 12 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 1 tconnect 1
<< end >>
