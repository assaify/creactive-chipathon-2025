** sch_path: /foss/designs/creactive-chipathon-2025/designs/libs/core_switch_matrix/switch_cell/switch_cell.sch
.subckt switch_cell DATA_IN CLK_PH1 CLK_PH2 EN DATA_OUT T1 T2 VDDD VSSD
*.PININFO DATA_IN:I CLK_PH1:I CLK_PH2:I DATA_OUT:O VDDD:B VSSD:B EN:I T1:B T2:B
x1 DATA_IN CLK_PH1 CLK_PH2 DATA_OUT VDDD VSSD dff_2ph_clk
x2 DATA_OUT EN VDDD VSSD T1 T2 tgate
.ends

* expanding   symbol:  libs/core_switch_matrix/dff_2ph_clk/dff_2ph_clk.sym # of pins=6
** sym_path: /foss/designs/creactive-chipathon-2025/designs/libs/core_switch_matrix/dff_2ph_clk/dff_2ph_clk.sym
** sch_path: /foss/designs/creactive-chipathon-2025/designs/libs/core_switch_matrix/dff_2ph_clk/dff_2ph_clk.sch
.subckt dff_2ph_clk D CLK_PH1 CLK_PH2 Q VDDD VSSD
*.PININFO D:I CLK_PH1:I CLK_PH2:I Q:O VDDD:B VSSD:B
x1 D CLK_PH1 net1 VDDD VDDD VSSD VSSD gf180mcu_fd_sc_mcu9t5v0__latq_1
x2 net1 CLK_PH2 Q VDDD VDDD VSSD VSSD gf180mcu_fd_sc_mcu9t5v0__latq_1
**** begin user architecture code

.include /foss/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/spice/gf180mcu_fd_sc_mcu9t5v0.spice

**** end user architecture code
.ends


* expanding   symbol:  libs/core_switch_matrix/tgate/tgate.sym # of pins=6
** sym_path: /foss/designs/creactive-chipathon-2025/designs/libs/core_switch_matrix/tgate/tgate.sym
** sch_path: /foss/designs/creactive-chipathon-2025/designs/libs/core_switch_matrix/tgate/tgate.sch
.subckt tgate CON EN VDDD VSSD T1 T2
*.PININFO CON:I EN:I VDDD:B VSSD:B T1:B T2:B
XM1 T2 NCON T1 VSSD nfet_03v3 L=0.28u W=4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=6
XM2 T2 PCON T1 VDDD pfet_03v3 L=0.28u W=4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=18
x1 CON EN net1 VDDD VDDD VSSD VSSD gf180mcu_fd_sc_mcu9t5v0__nand2_1
x2 net1 NCON VDDD VDDD VSSD VSSD gf180mcu_fd_sc_mcu9t5v0__inv_1
x3 NCON PCON VDDD VDDD VSSD VSSD gf180mcu_fd_sc_mcu9t5v0__inv_1
**** begin user architecture code

.include /foss/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu9t5v0/spice/gf180mcu_fd_sc_mcu9t5v0.spice

**** end user architecture code
.ends

