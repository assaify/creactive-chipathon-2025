magic
tech gf180mcuD
magscale 1 10
timestamp 1757672677
<< nwell >>
rect -352 -362 3204 1086
<< pmos >>
rect 38 0 94 800
rect 198 0 254 800
rect 358 0 414 800
rect 518 0 574 800
rect 678 0 734 800
rect 838 0 894 800
rect 998 0 1054 800
rect 1158 0 1214 800
rect 1318 0 1374 800
rect 1478 0 1534 800
rect 1638 0 1694 800
rect 1798 0 1854 800
rect 1958 0 2014 800
rect 2118 0 2174 800
rect 2278 0 2334 800
rect 2438 0 2494 800
rect 2598 0 2654 800
rect 2758 0 2814 800
<< pdiff >>
rect -92 729 38 800
rect -92 71 -69 729
rect -23 71 38 729
rect -92 0 38 71
rect 94 729 198 800
rect 94 71 123 729
rect 169 71 198 729
rect 94 0 198 71
rect 254 729 358 800
rect 254 71 283 729
rect 329 71 358 729
rect 254 0 358 71
rect 414 729 518 800
rect 414 71 443 729
rect 489 71 518 729
rect 414 0 518 71
rect 574 729 678 800
rect 574 71 603 729
rect 649 71 678 729
rect 574 0 678 71
rect 734 729 838 800
rect 734 71 763 729
rect 809 71 838 729
rect 734 0 838 71
rect 894 729 998 800
rect 894 71 923 729
rect 969 71 998 729
rect 894 0 998 71
rect 1054 729 1158 800
rect 1054 71 1083 729
rect 1129 71 1158 729
rect 1054 0 1158 71
rect 1214 729 1318 800
rect 1214 71 1243 729
rect 1289 71 1318 729
rect 1214 0 1318 71
rect 1374 729 1478 800
rect 1374 71 1403 729
rect 1449 71 1478 729
rect 1374 0 1478 71
rect 1534 729 1638 800
rect 1534 71 1563 729
rect 1609 71 1638 729
rect 1534 0 1638 71
rect 1694 729 1798 800
rect 1694 71 1723 729
rect 1769 71 1798 729
rect 1694 0 1798 71
rect 1854 729 1958 800
rect 1854 71 1883 729
rect 1929 71 1958 729
rect 1854 0 1958 71
rect 2014 729 2118 800
rect 2014 71 2043 729
rect 2089 71 2118 729
rect 2014 0 2118 71
rect 2174 729 2278 800
rect 2174 71 2203 729
rect 2249 71 2278 729
rect 2174 0 2278 71
rect 2334 729 2438 800
rect 2334 71 2363 729
rect 2409 71 2438 729
rect 2334 0 2438 71
rect 2494 729 2598 800
rect 2494 71 2523 729
rect 2569 71 2598 729
rect 2494 0 2598 71
rect 2654 729 2758 800
rect 2654 71 2683 729
rect 2729 71 2758 729
rect 2654 0 2758 71
rect 2814 729 2944 800
rect 2814 71 2875 729
rect 2921 71 2944 729
rect 2814 0 2944 71
<< pdiffc >>
rect -69 71 -23 729
rect 123 71 169 729
rect 283 71 329 729
rect 443 71 489 729
rect 603 71 649 729
rect 763 71 809 729
rect 923 71 969 729
rect 1083 71 1129 729
rect 1243 71 1289 729
rect 1403 71 1449 729
rect 1563 71 1609 729
rect 1723 71 1769 729
rect 1883 71 1929 729
rect 2043 71 2089 729
rect 2203 71 2249 729
rect 2363 71 2409 729
rect 2523 71 2569 729
rect 2683 71 2729 729
rect 2875 71 2921 729
<< nsubdiff >>
rect -264 983 3116 998
rect -264 937 -76 983
rect 2928 937 3116 983
rect -264 922 3116 937
rect -264 844 -188 922
rect -264 -120 -249 844
rect -203 -120 -188 844
rect 3040 844 3116 922
rect -264 -198 -188 -120
rect 3040 -120 3055 844
rect 3101 -120 3116 844
rect 3040 -198 3116 -120
rect -264 -213 3116 -198
rect -264 -259 -76 -213
rect 2928 -259 3116 -213
rect -264 -274 3116 -259
<< nsubdiffcont >>
rect -76 937 2928 983
rect -249 -120 -203 844
rect 3055 -120 3101 844
rect -76 -259 2928 -213
<< polysilicon >>
rect 38 800 94 860
rect 198 800 254 860
rect 358 800 414 860
rect 518 800 574 860
rect 678 800 734 860
rect 838 800 894 860
rect 998 800 1054 860
rect 1158 800 1214 860
rect 1318 800 1374 860
rect 1478 800 1534 860
rect 1638 800 1694 860
rect 1798 800 1854 860
rect 1958 800 2014 860
rect 2118 800 2174 860
rect 2278 800 2334 860
rect 2438 800 2494 860
rect 2598 800 2654 860
rect 2758 800 2814 860
rect 38 -60 94 0
rect 198 -60 254 0
rect 358 -60 414 0
rect 518 -60 574 0
rect 678 -60 734 0
rect 838 -60 894 0
rect 998 -60 1054 0
rect 1158 -60 1214 0
rect 1318 -60 1374 0
rect 1478 -60 1534 0
rect 1638 -60 1694 0
rect 1798 -60 1854 0
rect 1958 -60 2014 0
rect 2118 -60 2174 0
rect 2278 -60 2334 0
rect 2438 -60 2494 0
rect 2598 -60 2654 0
rect 2758 -60 2814 0
rect 28 -75 104 -60
rect 28 -121 43 -75
rect 89 -121 104 -75
rect 28 -136 104 -121
rect 188 -75 264 -60
rect 188 -121 203 -75
rect 249 -121 264 -75
rect 188 -136 264 -121
rect 348 -75 424 -60
rect 348 -121 363 -75
rect 409 -121 424 -75
rect 348 -136 424 -121
rect 508 -75 584 -60
rect 508 -121 523 -75
rect 569 -121 584 -75
rect 508 -136 584 -121
rect 668 -75 744 -60
rect 668 -121 683 -75
rect 729 -121 744 -75
rect 668 -136 744 -121
rect 828 -75 904 -60
rect 828 -121 843 -75
rect 889 -121 904 -75
rect 828 -136 904 -121
rect 988 -75 1064 -60
rect 988 -121 1003 -75
rect 1049 -121 1064 -75
rect 988 -136 1064 -121
rect 1148 -75 1224 -60
rect 1148 -121 1163 -75
rect 1209 -121 1224 -75
rect 1148 -136 1224 -121
rect 1308 -75 1384 -60
rect 1308 -121 1323 -75
rect 1369 -121 1384 -75
rect 1308 -136 1384 -121
rect 1468 -75 1544 -60
rect 1468 -121 1483 -75
rect 1529 -121 1544 -75
rect 1468 -136 1544 -121
rect 1628 -75 1704 -60
rect 1628 -121 1643 -75
rect 1689 -121 1704 -75
rect 1628 -136 1704 -121
rect 1788 -75 1864 -60
rect 1788 -121 1803 -75
rect 1849 -121 1864 -75
rect 1788 -136 1864 -121
rect 1948 -75 2024 -60
rect 1948 -121 1963 -75
rect 2009 -121 2024 -75
rect 1948 -136 2024 -121
rect 2108 -75 2184 -60
rect 2108 -121 2123 -75
rect 2169 -121 2184 -75
rect 2108 -136 2184 -121
rect 2268 -75 2344 -60
rect 2268 -121 2283 -75
rect 2329 -121 2344 -75
rect 2268 -136 2344 -121
rect 2428 -75 2504 -60
rect 2428 -121 2443 -75
rect 2489 -121 2504 -75
rect 2428 -136 2504 -121
rect 2588 -75 2664 -60
rect 2588 -121 2603 -75
rect 2649 -121 2664 -75
rect 2588 -136 2664 -121
rect 2748 -75 2824 -60
rect 2748 -121 2763 -75
rect 2809 -121 2824 -75
rect 2748 -136 2824 -121
<< polycontact >>
rect 43 -121 89 -75
rect 203 -121 249 -75
rect 363 -121 409 -75
rect 523 -121 569 -75
rect 683 -121 729 -75
rect 843 -121 889 -75
rect 1003 -121 1049 -75
rect 1163 -121 1209 -75
rect 1323 -121 1369 -75
rect 1483 -121 1529 -75
rect 1643 -121 1689 -75
rect 1803 -121 1849 -75
rect 1963 -121 2009 -75
rect 2123 -121 2169 -75
rect 2283 -121 2329 -75
rect 2443 -121 2489 -75
rect 2603 -121 2649 -75
rect 2763 -121 2809 -75
<< metal1 >>
rect -276 983 3128 1010
rect -276 937 -76 983
rect 2928 937 3128 983
rect -276 910 3128 937
rect -276 844 -176 910
rect -276 -120 -249 844
rect -203 -120 -176 844
rect 3028 844 3128 910
rect -84 729 -8 744
rect -84 71 -69 729
rect -23 71 -8 729
rect -84 56 -8 71
rect 108 729 184 744
rect 108 71 123 729
rect 169 71 184 729
rect 108 56 184 71
rect 268 729 344 744
rect 268 71 283 729
rect 329 71 344 729
rect 268 56 344 71
rect 428 729 504 744
rect 428 71 443 729
rect 489 71 504 729
rect 428 56 504 71
rect 588 729 664 744
rect 588 71 603 729
rect 649 71 664 729
rect 588 56 664 71
rect 748 729 824 744
rect 748 71 763 729
rect 809 71 824 729
rect 748 56 824 71
rect 908 729 984 744
rect 908 71 923 729
rect 969 71 984 729
rect 908 56 984 71
rect 1068 729 1144 744
rect 1068 71 1083 729
rect 1129 71 1144 729
rect 1068 56 1144 71
rect 1228 729 1304 744
rect 1228 71 1243 729
rect 1289 71 1304 729
rect 1228 56 1304 71
rect 1388 729 1464 744
rect 1388 71 1403 729
rect 1449 71 1464 729
rect 1388 56 1464 71
rect 1548 729 1624 744
rect 1548 71 1563 729
rect 1609 71 1624 729
rect 1548 56 1624 71
rect 1708 729 1784 744
rect 1708 71 1723 729
rect 1769 71 1784 729
rect 1708 56 1784 71
rect 1868 729 1944 744
rect 1868 71 1883 729
rect 1929 71 1944 729
rect 1868 56 1944 71
rect 2028 729 2104 744
rect 2028 71 2043 729
rect 2089 71 2104 729
rect 2028 56 2104 71
rect 2188 729 2264 744
rect 2188 71 2203 729
rect 2249 71 2264 729
rect 2188 56 2264 71
rect 2348 729 2424 744
rect 2348 71 2363 729
rect 2409 71 2424 729
rect 2348 56 2424 71
rect 2508 729 2584 744
rect 2508 71 2523 729
rect 2569 71 2584 729
rect 2508 56 2584 71
rect 2668 729 2744 744
rect 2668 71 2683 729
rect 2729 71 2744 729
rect 2668 56 2744 71
rect 2860 729 2936 744
rect 2860 71 2875 729
rect 2921 71 2936 729
rect 2860 56 2936 71
rect -276 -186 -176 -120
rect 28 -75 2824 -60
rect 28 -121 43 -75
rect 89 -121 203 -75
rect 249 -121 363 -75
rect 409 -121 523 -75
rect 569 -121 683 -75
rect 729 -121 843 -75
rect 889 -121 1003 -75
rect 1049 -121 1163 -75
rect 1209 -121 1323 -75
rect 1369 -121 1483 -75
rect 1529 -121 1643 -75
rect 1689 -121 1803 -75
rect 1849 -121 1963 -75
rect 2009 -121 2123 -75
rect 2169 -121 2283 -75
rect 2329 -121 2443 -75
rect 2489 -121 2603 -75
rect 2649 -121 2763 -75
rect 2809 -121 2824 -75
rect 28 -136 2824 -121
rect 3028 -120 3055 844
rect 3101 -120 3128 844
rect 3028 -186 3128 -120
rect -276 -213 3128 -186
rect -276 -259 -76 -213
rect 2928 -259 3128 -213
rect -276 -286 3128 -259
<< labels >>
flabel metal1 s 44 -120 44 -120 2 FreeSans 73 0 0 0 G
port 1 nsew
flabel metal1 s -68 72 -68 72 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 2876 72 2876 72 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 2524 72 2524 72 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 2204 72 2204 72 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 1884 72 1884 72 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 1564 73 1564 73 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 1244 73 1244 73 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 924 72 924 72 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 604 72 604 72 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 284 73 284 73 2 FreeSans 73 0 0 0 S
port 2 nsew
flabel metal1 s 2044 71 2044 71 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s 1724 71 1724 71 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s 1404 72 1404 72 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s 1084 72 1084 72 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s 764 71 764 71 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s 444 71 444 71 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s 124 72 124 72 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s 2364 71 2364 71 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s 2684 72 2684 72 2 FreeSans 73 0 0 0 D
port 3 nsew
flabel metal1 s -226 -236 -226 -236 2 FreeSans 73 0 0 0 B
port 4 nsew
<< properties >>
string path -1.490 4.800 15.390 4.800 15.390 -1.180 -1.130 -1.180 -1.130 4.440 
<< end >>
