magic
tech gf180mcuD
magscale 1 10
timestamp 1755277289
<< nwell >>
rect -1718 -4410 1718 4410
<< pmos >>
rect -1468 -4200 -1268 4200
rect -1164 -4200 -964 4200
rect -860 -4200 -660 4200
rect -556 -4200 -356 4200
rect -252 -4200 -52 4200
rect 52 -4200 252 4200
rect 356 -4200 556 4200
rect 660 -4200 860 4200
rect 964 -4200 1164 4200
rect 1268 -4200 1468 4200
<< pdiff >>
rect -1556 4187 -1468 4200
rect -1556 -4187 -1543 4187
rect -1497 -4187 -1468 4187
rect -1556 -4200 -1468 -4187
rect -1268 4187 -1164 4200
rect -1268 -4187 -1239 4187
rect -1193 -4187 -1164 4187
rect -1268 -4200 -1164 -4187
rect -964 4187 -860 4200
rect -964 -4187 -935 4187
rect -889 -4187 -860 4187
rect -964 -4200 -860 -4187
rect -660 4187 -556 4200
rect -660 -4187 -631 4187
rect -585 -4187 -556 4187
rect -660 -4200 -556 -4187
rect -356 4187 -252 4200
rect -356 -4187 -327 4187
rect -281 -4187 -252 4187
rect -356 -4200 -252 -4187
rect -52 4187 52 4200
rect -52 -4187 -23 4187
rect 23 -4187 52 4187
rect -52 -4200 52 -4187
rect 252 4187 356 4200
rect 252 -4187 281 4187
rect 327 -4187 356 4187
rect 252 -4200 356 -4187
rect 556 4187 660 4200
rect 556 -4187 585 4187
rect 631 -4187 660 4187
rect 556 -4200 660 -4187
rect 860 4187 964 4200
rect 860 -4187 889 4187
rect 935 -4187 964 4187
rect 860 -4200 964 -4187
rect 1164 4187 1268 4200
rect 1164 -4187 1193 4187
rect 1239 -4187 1268 4187
rect 1164 -4200 1268 -4187
rect 1468 4187 1556 4200
rect 1468 -4187 1497 4187
rect 1543 -4187 1556 4187
rect 1468 -4200 1556 -4187
<< pdiffc >>
rect -1543 -4187 -1497 4187
rect -1239 -4187 -1193 4187
rect -935 -4187 -889 4187
rect -631 -4187 -585 4187
rect -327 -4187 -281 4187
rect -23 -4187 23 4187
rect 281 -4187 327 4187
rect 585 -4187 631 4187
rect 889 -4187 935 4187
rect 1193 -4187 1239 4187
rect 1497 -4187 1543 4187
<< nsubdiff >>
rect -1694 4314 1694 4386
rect -1694 4270 -1622 4314
rect -1694 -4270 -1681 4270
rect -1635 -4270 -1622 4270
rect 1622 4270 1694 4314
rect -1694 -4314 -1622 -4270
rect 1622 -4270 1635 4270
rect 1681 -4270 1694 4270
rect 1622 -4314 1694 -4270
rect -1694 -4386 1694 -4314
<< nsubdiffcont >>
rect -1681 -4270 -1635 4270
rect 1635 -4270 1681 4270
<< polysilicon >>
rect -1468 4279 -1268 4292
rect -1468 4233 -1455 4279
rect -1281 4233 -1268 4279
rect -1468 4200 -1268 4233
rect -1164 4279 -964 4292
rect -1164 4233 -1151 4279
rect -977 4233 -964 4279
rect -1164 4200 -964 4233
rect -860 4279 -660 4292
rect -860 4233 -847 4279
rect -673 4233 -660 4279
rect -860 4200 -660 4233
rect -556 4279 -356 4292
rect -556 4233 -543 4279
rect -369 4233 -356 4279
rect -556 4200 -356 4233
rect -252 4279 -52 4292
rect -252 4233 -239 4279
rect -65 4233 -52 4279
rect -252 4200 -52 4233
rect 52 4279 252 4292
rect 52 4233 65 4279
rect 239 4233 252 4279
rect 52 4200 252 4233
rect 356 4279 556 4292
rect 356 4233 369 4279
rect 543 4233 556 4279
rect 356 4200 556 4233
rect 660 4279 860 4292
rect 660 4233 673 4279
rect 847 4233 860 4279
rect 660 4200 860 4233
rect 964 4279 1164 4292
rect 964 4233 977 4279
rect 1151 4233 1164 4279
rect 964 4200 1164 4233
rect 1268 4279 1468 4292
rect 1268 4233 1281 4279
rect 1455 4233 1468 4279
rect 1268 4200 1468 4233
rect -1468 -4233 -1268 -4200
rect -1468 -4279 -1455 -4233
rect -1281 -4279 -1268 -4233
rect -1468 -4292 -1268 -4279
rect -1164 -4233 -964 -4200
rect -1164 -4279 -1151 -4233
rect -977 -4279 -964 -4233
rect -1164 -4292 -964 -4279
rect -860 -4233 -660 -4200
rect -860 -4279 -847 -4233
rect -673 -4279 -660 -4233
rect -860 -4292 -660 -4279
rect -556 -4233 -356 -4200
rect -556 -4279 -543 -4233
rect -369 -4279 -356 -4233
rect -556 -4292 -356 -4279
rect -252 -4233 -52 -4200
rect -252 -4279 -239 -4233
rect -65 -4279 -52 -4233
rect -252 -4292 -52 -4279
rect 52 -4233 252 -4200
rect 52 -4279 65 -4233
rect 239 -4279 252 -4233
rect 52 -4292 252 -4279
rect 356 -4233 556 -4200
rect 356 -4279 369 -4233
rect 543 -4279 556 -4233
rect 356 -4292 556 -4279
rect 660 -4233 860 -4200
rect 660 -4279 673 -4233
rect 847 -4279 860 -4233
rect 660 -4292 860 -4279
rect 964 -4233 1164 -4200
rect 964 -4279 977 -4233
rect 1151 -4279 1164 -4233
rect 964 -4292 1164 -4279
rect 1268 -4233 1468 -4200
rect 1268 -4279 1281 -4233
rect 1455 -4279 1468 -4233
rect 1268 -4292 1468 -4279
<< polycontact >>
rect -1455 4233 -1281 4279
rect -1151 4233 -977 4279
rect -847 4233 -673 4279
rect -543 4233 -369 4279
rect -239 4233 -65 4279
rect 65 4233 239 4279
rect 369 4233 543 4279
rect 673 4233 847 4279
rect 977 4233 1151 4279
rect 1281 4233 1455 4279
rect -1455 -4279 -1281 -4233
rect -1151 -4279 -977 -4233
rect -847 -4279 -673 -4233
rect -543 -4279 -369 -4233
rect -239 -4279 -65 -4233
rect 65 -4279 239 -4233
rect 369 -4279 543 -4233
rect 673 -4279 847 -4233
rect 977 -4279 1151 -4233
rect 1281 -4279 1455 -4233
<< metal1 >>
rect -1681 4327 1681 4373
rect -1681 4270 -1635 4327
rect -1466 4233 -1455 4279
rect -1281 4233 -1270 4279
rect -1162 4233 -1151 4279
rect -977 4233 -966 4279
rect -858 4233 -847 4279
rect -673 4233 -662 4279
rect -554 4233 -543 4279
rect -369 4233 -358 4279
rect -250 4233 -239 4279
rect -65 4233 -54 4279
rect 54 4233 65 4279
rect 239 4233 250 4279
rect 358 4233 369 4279
rect 543 4233 554 4279
rect 662 4233 673 4279
rect 847 4233 858 4279
rect 966 4233 977 4279
rect 1151 4233 1162 4279
rect 1270 4233 1281 4279
rect 1455 4233 1466 4279
rect 1635 4270 1681 4327
rect -1543 4187 -1497 4198
rect -1543 -4198 -1497 -4187
rect -1239 4187 -1193 4198
rect -1239 -4198 -1193 -4187
rect -935 4187 -889 4198
rect -935 -4198 -889 -4187
rect -631 4187 -585 4198
rect -631 -4198 -585 -4187
rect -327 4187 -281 4198
rect -327 -4198 -281 -4187
rect -23 4187 23 4198
rect -23 -4198 23 -4187
rect 281 4187 327 4198
rect 281 -4198 327 -4187
rect 585 4187 631 4198
rect 585 -4198 631 -4187
rect 889 4187 935 4198
rect 889 -4198 935 -4187
rect 1193 4187 1239 4198
rect 1193 -4198 1239 -4187
rect 1497 4187 1543 4198
rect 1497 -4198 1543 -4187
rect -1681 -4327 -1635 -4270
rect -1466 -4279 -1455 -4233
rect -1281 -4279 -1270 -4233
rect -1162 -4279 -1151 -4233
rect -977 -4279 -966 -4233
rect -858 -4279 -847 -4233
rect -673 -4279 -662 -4233
rect -554 -4279 -543 -4233
rect -369 -4279 -358 -4233
rect -250 -4279 -239 -4233
rect -65 -4279 -54 -4233
rect 54 -4279 65 -4233
rect 239 -4279 250 -4233
rect 358 -4279 369 -4233
rect 543 -4279 554 -4233
rect 662 -4279 673 -4233
rect 847 -4279 858 -4233
rect 966 -4279 977 -4233
rect 1151 -4279 1162 -4233
rect 1270 -4279 1281 -4233
rect 1455 -4279 1466 -4233
rect 1635 -4327 1681 -4270
rect -1681 -4373 1681 -4327
<< properties >>
string FIXED_BBOX -1658 -4350 1658 4350
string gencell pfet_03v3
string library gf180mcu
string parameters w 42.0 l 1.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0}
<< end >>
