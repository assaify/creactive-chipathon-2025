magic
tech gf180mcuD
magscale 1 10
timestamp 1755277289
<< pwell >>
rect -806 -435 806 435
<< nmos >>
rect -556 -225 -356 225
rect -252 -225 -52 225
rect 52 -225 252 225
rect 356 -225 556 225
<< ndiff >>
rect -644 212 -556 225
rect -644 -212 -631 212
rect -585 -212 -556 212
rect -644 -225 -556 -212
rect -356 212 -252 225
rect -356 -212 -327 212
rect -281 -212 -252 212
rect -356 -225 -252 -212
rect -52 212 52 225
rect -52 -212 -23 212
rect 23 -212 52 212
rect -52 -225 52 -212
rect 252 212 356 225
rect 252 -212 281 212
rect 327 -212 356 212
rect 252 -225 356 -212
rect 556 212 644 225
rect 556 -212 585 212
rect 631 -212 644 212
rect 556 -225 644 -212
<< ndiffc >>
rect -631 -212 -585 212
rect -327 -212 -281 212
rect -23 -212 23 212
rect 281 -212 327 212
rect 585 -212 631 212
<< psubdiff >>
rect -782 339 782 411
rect -782 295 -710 339
rect -782 -295 -769 295
rect -723 -295 -710 295
rect 710 295 782 339
rect -782 -339 -710 -295
rect 710 -295 723 295
rect 769 -295 782 295
rect 710 -339 782 -295
rect -782 -411 782 -339
<< psubdiffcont >>
rect -769 -295 -723 295
rect 723 -295 769 295
<< polysilicon >>
rect -556 304 -356 317
rect -556 258 -543 304
rect -369 258 -356 304
rect -556 225 -356 258
rect -252 304 -52 317
rect -252 258 -239 304
rect -65 258 -52 304
rect -252 225 -52 258
rect 52 304 252 317
rect 52 258 65 304
rect 239 258 252 304
rect 52 225 252 258
rect 356 304 556 317
rect 356 258 369 304
rect 543 258 556 304
rect 356 225 556 258
rect -556 -258 -356 -225
rect -556 -304 -543 -258
rect -369 -304 -356 -258
rect -556 -317 -356 -304
rect -252 -258 -52 -225
rect -252 -304 -239 -258
rect -65 -304 -52 -258
rect -252 -317 -52 -304
rect 52 -258 252 -225
rect 52 -304 65 -258
rect 239 -304 252 -258
rect 52 -317 252 -304
rect 356 -258 556 -225
rect 356 -304 369 -258
rect 543 -304 556 -258
rect 356 -317 556 -304
<< polycontact >>
rect -543 258 -369 304
rect -239 258 -65 304
rect 65 258 239 304
rect 369 258 543 304
rect -543 -304 -369 -258
rect -239 -304 -65 -258
rect 65 -304 239 -258
rect 369 -304 543 -258
<< metal1 >>
rect -769 352 769 398
rect -769 295 -723 352
rect -554 258 -543 304
rect -369 258 -358 304
rect -250 258 -239 304
rect -65 258 -54 304
rect 54 258 65 304
rect 239 258 250 304
rect 358 258 369 304
rect 543 258 554 304
rect 723 295 769 352
rect -631 212 -585 223
rect -631 -223 -585 -212
rect -327 212 -281 223
rect -327 -223 -281 -212
rect -23 212 23 223
rect -23 -223 23 -212
rect 281 212 327 223
rect 281 -223 327 -212
rect 585 212 631 223
rect 585 -223 631 -212
rect -769 -352 -723 -295
rect -554 -304 -543 -258
rect -369 -304 -358 -258
rect -250 -304 -239 -258
rect -65 -304 -54 -258
rect 54 -304 65 -258
rect 239 -304 250 -258
rect 358 -304 369 -258
rect 543 -304 554 -258
rect 723 -352 769 -295
rect -769 -398 769 -352
<< properties >>
string FIXED_BBOX -746 -375 746 375
string gencell nfet_03v3
string library gf180mcu
string parameters w 2.25 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
