magic
tech gf180mcuD
magscale 1 10
timestamp 1755276408
<< nwell >>
rect -350 -43254 350 43254
<< pmos >>
rect -100 34644 100 43044
rect -100 26012 100 34412
rect -100 17380 100 25780
rect -100 8748 100 17148
rect -100 116 100 8516
rect -100 -8516 100 -116
rect -100 -17148 100 -8748
rect -100 -25780 100 -17380
rect -100 -34412 100 -26012
rect -100 -43044 100 -34644
<< pdiff >>
rect -188 43031 -100 43044
rect -188 34657 -175 43031
rect -129 34657 -100 43031
rect -188 34644 -100 34657
rect 100 43031 188 43044
rect 100 34657 129 43031
rect 175 34657 188 43031
rect 100 34644 188 34657
rect -188 34399 -100 34412
rect -188 26025 -175 34399
rect -129 26025 -100 34399
rect -188 26012 -100 26025
rect 100 34399 188 34412
rect 100 26025 129 34399
rect 175 26025 188 34399
rect 100 26012 188 26025
rect -188 25767 -100 25780
rect -188 17393 -175 25767
rect -129 17393 -100 25767
rect -188 17380 -100 17393
rect 100 25767 188 25780
rect 100 17393 129 25767
rect 175 17393 188 25767
rect 100 17380 188 17393
rect -188 17135 -100 17148
rect -188 8761 -175 17135
rect -129 8761 -100 17135
rect -188 8748 -100 8761
rect 100 17135 188 17148
rect 100 8761 129 17135
rect 175 8761 188 17135
rect 100 8748 188 8761
rect -188 8503 -100 8516
rect -188 129 -175 8503
rect -129 129 -100 8503
rect -188 116 -100 129
rect 100 8503 188 8516
rect 100 129 129 8503
rect 175 129 188 8503
rect 100 116 188 129
rect -188 -129 -100 -116
rect -188 -8503 -175 -129
rect -129 -8503 -100 -129
rect -188 -8516 -100 -8503
rect 100 -129 188 -116
rect 100 -8503 129 -129
rect 175 -8503 188 -129
rect 100 -8516 188 -8503
rect -188 -8761 -100 -8748
rect -188 -17135 -175 -8761
rect -129 -17135 -100 -8761
rect -188 -17148 -100 -17135
rect 100 -8761 188 -8748
rect 100 -17135 129 -8761
rect 175 -17135 188 -8761
rect 100 -17148 188 -17135
rect -188 -17393 -100 -17380
rect -188 -25767 -175 -17393
rect -129 -25767 -100 -17393
rect -188 -25780 -100 -25767
rect 100 -17393 188 -17380
rect 100 -25767 129 -17393
rect 175 -25767 188 -17393
rect 100 -25780 188 -25767
rect -188 -26025 -100 -26012
rect -188 -34399 -175 -26025
rect -129 -34399 -100 -26025
rect -188 -34412 -100 -34399
rect 100 -26025 188 -26012
rect 100 -34399 129 -26025
rect 175 -34399 188 -26025
rect 100 -34412 188 -34399
rect -188 -34657 -100 -34644
rect -188 -43031 -175 -34657
rect -129 -43031 -100 -34657
rect -188 -43044 -100 -43031
rect 100 -34657 188 -34644
rect 100 -43031 129 -34657
rect 175 -43031 188 -34657
rect 100 -43044 188 -43031
<< pdiffc >>
rect -175 34657 -129 43031
rect 129 34657 175 43031
rect -175 26025 -129 34399
rect 129 26025 175 34399
rect -175 17393 -129 25767
rect 129 17393 175 25767
rect -175 8761 -129 17135
rect 129 8761 175 17135
rect -175 129 -129 8503
rect 129 129 175 8503
rect -175 -8503 -129 -129
rect 129 -8503 175 -129
rect -175 -17135 -129 -8761
rect 129 -17135 175 -8761
rect -175 -25767 -129 -17393
rect 129 -25767 175 -17393
rect -175 -34399 -129 -26025
rect 129 -34399 175 -26025
rect -175 -43031 -129 -34657
rect 129 -43031 175 -34657
<< nsubdiff >>
rect -326 43158 326 43230
rect -326 43114 -254 43158
rect -326 -43114 -313 43114
rect -267 -43114 -254 43114
rect 254 43114 326 43158
rect -326 -43158 -254 -43114
rect 254 -43114 267 43114
rect 313 -43114 326 43114
rect 254 -43158 326 -43114
rect -326 -43230 326 -43158
<< nsubdiffcont >>
rect -313 -43114 -267 43114
rect 267 -43114 313 43114
<< polysilicon >>
rect -100 43123 100 43136
rect -100 43077 -87 43123
rect 87 43077 100 43123
rect -100 43044 100 43077
rect -100 34611 100 34644
rect -100 34565 -87 34611
rect 87 34565 100 34611
rect -100 34552 100 34565
rect -100 34491 100 34504
rect -100 34445 -87 34491
rect 87 34445 100 34491
rect -100 34412 100 34445
rect -100 25979 100 26012
rect -100 25933 -87 25979
rect 87 25933 100 25979
rect -100 25920 100 25933
rect -100 25859 100 25872
rect -100 25813 -87 25859
rect 87 25813 100 25859
rect -100 25780 100 25813
rect -100 17347 100 17380
rect -100 17301 -87 17347
rect 87 17301 100 17347
rect -100 17288 100 17301
rect -100 17227 100 17240
rect -100 17181 -87 17227
rect 87 17181 100 17227
rect -100 17148 100 17181
rect -100 8715 100 8748
rect -100 8669 -87 8715
rect 87 8669 100 8715
rect -100 8656 100 8669
rect -100 8595 100 8608
rect -100 8549 -87 8595
rect 87 8549 100 8595
rect -100 8516 100 8549
rect -100 83 100 116
rect -100 37 -87 83
rect 87 37 100 83
rect -100 24 100 37
rect -100 -37 100 -24
rect -100 -83 -87 -37
rect 87 -83 100 -37
rect -100 -116 100 -83
rect -100 -8549 100 -8516
rect -100 -8595 -87 -8549
rect 87 -8595 100 -8549
rect -100 -8608 100 -8595
rect -100 -8669 100 -8656
rect -100 -8715 -87 -8669
rect 87 -8715 100 -8669
rect -100 -8748 100 -8715
rect -100 -17181 100 -17148
rect -100 -17227 -87 -17181
rect 87 -17227 100 -17181
rect -100 -17240 100 -17227
rect -100 -17301 100 -17288
rect -100 -17347 -87 -17301
rect 87 -17347 100 -17301
rect -100 -17380 100 -17347
rect -100 -25813 100 -25780
rect -100 -25859 -87 -25813
rect 87 -25859 100 -25813
rect -100 -25872 100 -25859
rect -100 -25933 100 -25920
rect -100 -25979 -87 -25933
rect 87 -25979 100 -25933
rect -100 -26012 100 -25979
rect -100 -34445 100 -34412
rect -100 -34491 -87 -34445
rect 87 -34491 100 -34445
rect -100 -34504 100 -34491
rect -100 -34565 100 -34552
rect -100 -34611 -87 -34565
rect 87 -34611 100 -34565
rect -100 -34644 100 -34611
rect -100 -43077 100 -43044
rect -100 -43123 -87 -43077
rect 87 -43123 100 -43077
rect -100 -43136 100 -43123
<< polycontact >>
rect -87 43077 87 43123
rect -87 34565 87 34611
rect -87 34445 87 34491
rect -87 25933 87 25979
rect -87 25813 87 25859
rect -87 17301 87 17347
rect -87 17181 87 17227
rect -87 8669 87 8715
rect -87 8549 87 8595
rect -87 37 87 83
rect -87 -83 87 -37
rect -87 -8595 87 -8549
rect -87 -8715 87 -8669
rect -87 -17227 87 -17181
rect -87 -17347 87 -17301
rect -87 -25859 87 -25813
rect -87 -25979 87 -25933
rect -87 -34491 87 -34445
rect -87 -34611 87 -34565
rect -87 -43123 87 -43077
<< metal1 >>
rect -313 43171 313 43217
rect -313 43114 -267 43171
rect -98 43077 -87 43123
rect 87 43077 98 43123
rect 267 43114 313 43171
rect -175 43031 -129 43042
rect -175 34646 -129 34657
rect 129 43031 175 43042
rect 129 34646 175 34657
rect -98 34565 -87 34611
rect 87 34565 98 34611
rect -98 34445 -87 34491
rect 87 34445 98 34491
rect -175 34399 -129 34410
rect -175 26014 -129 26025
rect 129 34399 175 34410
rect 129 26014 175 26025
rect -98 25933 -87 25979
rect 87 25933 98 25979
rect -98 25813 -87 25859
rect 87 25813 98 25859
rect -175 25767 -129 25778
rect -175 17382 -129 17393
rect 129 25767 175 25778
rect 129 17382 175 17393
rect -98 17301 -87 17347
rect 87 17301 98 17347
rect -98 17181 -87 17227
rect 87 17181 98 17227
rect -175 17135 -129 17146
rect -175 8750 -129 8761
rect 129 17135 175 17146
rect 129 8750 175 8761
rect -98 8669 -87 8715
rect 87 8669 98 8715
rect -98 8549 -87 8595
rect 87 8549 98 8595
rect -175 8503 -129 8514
rect -175 118 -129 129
rect 129 8503 175 8514
rect 129 118 175 129
rect -98 37 -87 83
rect 87 37 98 83
rect -98 -83 -87 -37
rect 87 -83 98 -37
rect -175 -129 -129 -118
rect -175 -8514 -129 -8503
rect 129 -129 175 -118
rect 129 -8514 175 -8503
rect -98 -8595 -87 -8549
rect 87 -8595 98 -8549
rect -98 -8715 -87 -8669
rect 87 -8715 98 -8669
rect -175 -8761 -129 -8750
rect -175 -17146 -129 -17135
rect 129 -8761 175 -8750
rect 129 -17146 175 -17135
rect -98 -17227 -87 -17181
rect 87 -17227 98 -17181
rect -98 -17347 -87 -17301
rect 87 -17347 98 -17301
rect -175 -17393 -129 -17382
rect -175 -25778 -129 -25767
rect 129 -17393 175 -17382
rect 129 -25778 175 -25767
rect -98 -25859 -87 -25813
rect 87 -25859 98 -25813
rect -98 -25979 -87 -25933
rect 87 -25979 98 -25933
rect -175 -26025 -129 -26014
rect -175 -34410 -129 -34399
rect 129 -26025 175 -26014
rect 129 -34410 175 -34399
rect -98 -34491 -87 -34445
rect 87 -34491 98 -34445
rect -98 -34611 -87 -34565
rect 87 -34611 98 -34565
rect -175 -34657 -129 -34646
rect -175 -43042 -129 -43031
rect 129 -34657 175 -34646
rect 129 -43042 175 -43031
rect -313 -43171 -267 -43114
rect -98 -43123 -87 -43077
rect 87 -43123 98 -43077
rect 267 -43171 313 -43114
rect -313 -43217 313 -43171
<< properties >>
string FIXED_BBOX -290 -43194 290 43194
string gencell pfet_03v3
string library gf180mcu
string parameters w 42.0 l 1.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
