magic
tech gf180mcuD
magscale 1 10
timestamp 1757676927
<< error_s >>
rect -322 1010 -284 1056
rect -276 998 -238 1010
rect -105 998 -67 1012
rect 1010 998 1066 1012
rect 1170 998 1226 1012
rect 1330 998 1386 1012
rect 1490 998 1546 1012
rect 1650 998 1706 1012
rect 1810 998 1866 1012
rect -276 983 1996 998
rect 2107 983 2153 1304
rect -276 937 2928 983
rect -276 922 2184 937
rect -276 893 -180 922
rect -276 531 -147 893
rect -25 800 0 922
rect 2 889 21 922
rect 56 918 370 922
rect 50 902 370 918
rect 426 902 504 922
rect 3 816 36 862
rect 37 849 517 902
rect 530 860 533 918
rect 615 862 661 922
rect 775 910 821 922
rect 518 849 533 860
rect 37 800 592 849
rect 600 800 661 862
rect 678 852 690 860
rect 697 852 722 910
rect 760 896 821 910
rect 760 852 850 896
rect 920 852 1010 922
rect 1112 874 1188 922
rect 1112 852 1202 874
rect 1240 852 1246 910
rect 1255 852 1301 922
rect 1415 896 1461 922
rect 1575 910 1621 922
rect 1318 852 1330 860
rect 1386 852 1464 896
rect 1478 852 1490 860
rect 1493 852 1522 910
rect 1560 896 1621 910
rect 1560 852 1650 896
rect 678 800 1781 852
rect -130 744 -124 790
rect -84 758 1781 800
rect -98 729 1781 758
rect -84 652 1781 729
rect -276 516 -180 531
rect -264 460 -180 516
rect -84 460 1026 652
rect 1049 636 1058 652
rect 1083 472 1202 652
rect 1214 608 1224 652
rect 1214 520 1223 608
rect 1243 576 1781 652
rect 1243 531 1301 576
rect 1318 531 1330 576
rect 1374 532 1464 576
rect 1243 472 1289 531
rect -264 304 -188 460
rect -256 262 -188 304
rect -180 262 -156 460
rect -92 453 1026 460
rect 1054 453 1202 472
rect 1214 453 1289 472
rect 1403 521 1464 532
rect 1478 531 1490 576
rect 1563 532 1650 576
rect 1563 531 1621 532
rect 1628 531 1650 532
rect 1723 531 1781 576
rect 1798 531 1810 860
rect 1908 800 2002 922
rect 2092 860 2168 922
rect 2092 800 2174 860
rect 1854 729 1866 758
rect 1883 574 1895 729
rect 1908 574 2184 800
rect 1883 573 2184 574
rect 1883 531 2002 573
rect 1403 516 1476 521
rect 1374 453 1386 460
rect 1403 453 1464 516
rect 1534 453 1546 460
rect 1563 453 1609 531
rect 1628 521 1638 531
rect 1624 516 1638 521
rect 1628 453 1638 516
rect 1723 465 1769 531
rect 1784 516 1796 519
rect 1868 465 1869 519
rect 1883 465 1929 531
rect 1694 453 1798 465
rect 1854 453 1958 465
rect 2014 453 2174 573
rect 2188 453 2226 744
rect -256 247 -180 262
rect -1024 206 -180 247
rect -1300 201 -180 206
rect -1300 98 -352 201
rect -256 186 -180 201
rect -256 -5 -188 186
rect -180 -5 -156 186
rect -92 0 2326 453
rect -256 -25 -156 -5
rect -256 -64 -166 -25
rect -991 -90 -747 -64
rect -701 -90 -276 -64
rect -256 -69 -115 -64
rect -264 -90 -115 -69
rect -86 -86 2326 0
rect -69 -90 28 -86
rect -264 -119 -166 -90
rect -264 -120 -174 -119
rect -264 -196 -180 -120
rect 43 -121 89 -86
rect 203 -121 249 -86
rect 363 -121 409 -86
rect 523 -121 569 -86
rect 683 -89 762 -86
rect 683 -121 777 -89
rect 716 -156 777 -121
rect 716 -172 717 -156
rect -56 -196 717 -172
rect -264 -198 -56 -196
rect 731 -198 777 -156
rect 792 -172 816 -86
rect 843 -121 889 -86
rect 904 -90 988 -86
rect 1010 -90 1127 -86
rect 904 -119 1127 -90
rect 1148 -90 1308 -86
rect 1330 -90 1468 -86
rect 1490 -90 1628 -86
rect 1650 -90 1788 -86
rect 1810 -90 1948 -86
rect 1148 -119 1948 -90
rect 904 -134 1948 -119
rect 888 -154 924 -134
rect 968 -136 1010 -134
rect 968 -154 988 -136
rect 888 -156 908 -154
rect 888 -172 889 -156
rect 792 -196 889 -172
rect 1010 -184 1028 -182
rect 1112 -184 1188 -134
rect 1288 -136 1330 -134
rect 1448 -136 1490 -134
rect 1608 -136 1650 -134
rect 1768 -136 1810 -134
rect 1928 -136 1988 -134
rect 1288 -154 1308 -136
rect 1448 -154 1468 -136
rect 1608 -154 1628 -136
rect 1768 -154 1788 -136
rect 1928 -154 1948 -136
rect 1968 -156 2074 -136
rect 1010 -196 1066 -184
rect 1112 -196 1226 -184
rect 888 -198 1226 -196
rect 1330 -198 1386 -184
rect 1490 -198 1546 -184
rect 1650 -198 1706 -184
rect 1810 -198 1866 -184
rect 1988 -198 2074 -156
rect 2084 -198 2085 -86
rect 2099 -89 2160 -86
rect 2108 -121 2160 -89
rect 2108 -136 2174 -121
rect 2140 -156 2184 -136
rect 2160 -198 2184 -156
rect -747 -262 -701 -203
rect -1169 -280 -1145 -271
rect -1016 -280 -946 -262
rect -1169 -290 -1121 -280
rect -1075 -290 -946 -280
rect -1169 -319 -1145 -290
rect -1121 -326 -1075 -290
rect -1016 -306 -946 -290
rect -776 -297 -701 -262
rect -264 -272 1988 -198
rect -264 -274 -55 -272
rect 72 -274 393 -272
rect 716 -274 792 -272
rect 888 -274 1988 -272
rect 2084 -274 2160 -198
rect -672 -297 -667 -290
rect -776 -306 -667 -297
rect -115 -299 -114 -274
rect -1121 -343 -1046 -326
rect -747 -343 -667 -306
rect -319 -343 -273 -299
rect -1116 -356 -1046 -343
rect -2037 -440 -2035 -430
rect -2035 -450 -2025 -440
rect -2039 -496 -2037 -494
rect -2035 -496 -2025 -486
rect -1134 -488 -1046 -356
rect -713 -365 -667 -343
rect -1043 -470 -1029 -372
rect -876 -476 -842 -424
rect -611 -432 -484 -365
rect -698 -476 -654 -432
rect -714 -487 -654 -476
rect -869 -488 -654 -487
rect -2039 -506 -2035 -496
rect -2039 -635 -2037 -506
rect -1134 -536 -1074 -488
rect -869 -533 -865 -488
rect -1134 -555 -1046 -536
rect -823 -555 -819 -533
rect -714 -536 -654 -488
rect -672 -555 -654 -536
rect -539 -476 -467 -437
rect -539 -483 -512 -476
rect -539 -543 -467 -483
rect -331 -487 -272 -483
rect -331 -496 -271 -487
rect -331 -543 -254 -496
rect -244 -543 -243 -318
rect -115 -343 -69 -299
rect 117 -523 144 -274
rect 716 -362 717 -274
rect 792 -362 816 -274
rect 888 -362 889 -274
rect 1988 -362 2074 -274
rect 2084 -362 2085 -274
rect 2160 -362 2184 -274
rect -539 -555 -451 -543
rect -331 -555 -243 -543
rect -1427 -742 -1425 -598
rect -1429 -752 -1425 -742
rect -1439 -762 -1429 -752
rect -1427 -754 -1425 -752
rect -1257 -755 310 -555
rect -916 -761 -836 -755
rect -1439 -808 -1429 -798
rect -976 -803 -836 -761
rect -386 -778 -184 -755
rect -591 -785 -553 -780
rect -661 -802 -613 -785
rect -1429 -818 -1427 -808
rect -976 -821 -886 -803
rect -976 -831 -946 -821
rect -842 -831 -836 -803
rect -507 -803 -423 -780
rect -386 -802 -371 -778
rect -507 -813 -404 -803
rect -976 -875 -926 -831
rect -862 -875 -836 -831
rect -555 -851 -492 -835
rect -555 -864 -467 -851
rect -687 -888 -641 -873
rect -1096 -945 -1046 -901
rect -742 -945 -716 -892
rect -539 -901 -467 -864
rect -423 -875 -404 -813
rect -306 -831 -254 -778
rect -230 -802 -184 -778
rect -174 -802 -150 -755
rect -245 -831 -184 -802
rect -306 -842 -184 -831
rect -306 -860 -208 -842
rect -263 -864 -208 -860
rect -319 -872 -208 -864
rect -263 -875 -244 -872
rect 125 -873 144 -771
rect -351 -901 -332 -875
rect -672 -1005 -654 -901
rect -539 -945 -492 -901
rect -143 -921 -124 -892
rect 85 -898 144 -873
rect -114 -939 -95 -921
rect 97 -926 144 -898
rect -539 -1005 -479 -945
rect -143 -983 -124 -939
rect -1270 -1098 -1121 -1072
rect -1075 -1098 -545 -1072
rect -469 -1098 -338 -1072
rect -292 -1098 110 -1072
rect 156 -1098 224 -1072
rect -1257 -1294 310 -1206
rect -2039 -1927 -2037 -1796
rect -256 -2152 -254 -1874
use dff_2ph_clk$1  dff_2ph_clk$1_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -2326 -2405 310 103
use gf180mcu_fd_sc_mcu9t5v0__fill_2  gf180mcu_fd_sc_mcu9t5v0__fill_2_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie$1  gf180mcu_fd_sc_mcu9t5v0__filltie$1_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__filltie  gf180mcu_fd_sc_mcu9t5v0__filltie_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  gf180mcu_fd_sc_mcu9t5v0__inv_1_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__latq_1  gf180mcu_fd_sc_mcu9t5v0__latq_1_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -86 -90 2326 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  gf180mcu_fd_sc_mcu9t5v0__nand2_1_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -86 -90 646 1098
use nfet  nfet_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -268 -284 1200 1010
use pfet  pfet_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -352 -362 3204 1086
use tgate$1  tgate$1_0
timestamp 1757676927
transform 1 0 0 0 1 0
box -1300 -1318 2256 1570
<< end >>
