magic
tech gf180mcuD
magscale 1 10
timestamp 1755276408
<< pwell >>
rect -350 -1458 350 1458
<< nmos >>
rect -100 798 100 1248
rect -100 116 100 566
rect -100 -566 100 -116
rect -100 -1248 100 -798
<< ndiff >>
rect -188 1235 -100 1248
rect -188 811 -175 1235
rect -129 811 -100 1235
rect -188 798 -100 811
rect 100 1235 188 1248
rect 100 811 129 1235
rect 175 811 188 1235
rect 100 798 188 811
rect -188 553 -100 566
rect -188 129 -175 553
rect -129 129 -100 553
rect -188 116 -100 129
rect 100 553 188 566
rect 100 129 129 553
rect 175 129 188 553
rect 100 116 188 129
rect -188 -129 -100 -116
rect -188 -553 -175 -129
rect -129 -553 -100 -129
rect -188 -566 -100 -553
rect 100 -129 188 -116
rect 100 -553 129 -129
rect 175 -553 188 -129
rect 100 -566 188 -553
rect -188 -811 -100 -798
rect -188 -1235 -175 -811
rect -129 -1235 -100 -811
rect -188 -1248 -100 -1235
rect 100 -811 188 -798
rect 100 -1235 129 -811
rect 175 -1235 188 -811
rect 100 -1248 188 -1235
<< ndiffc >>
rect -175 811 -129 1235
rect 129 811 175 1235
rect -175 129 -129 553
rect 129 129 175 553
rect -175 -553 -129 -129
rect 129 -553 175 -129
rect -175 -1235 -129 -811
rect 129 -1235 175 -811
<< psubdiff >>
rect -326 1362 326 1434
rect -326 1318 -254 1362
rect -326 -1318 -313 1318
rect -267 -1318 -254 1318
rect 254 1318 326 1362
rect -326 -1362 -254 -1318
rect 254 -1318 267 1318
rect 313 -1318 326 1318
rect 254 -1362 326 -1318
rect -326 -1434 326 -1362
<< psubdiffcont >>
rect -313 -1318 -267 1318
rect 267 -1318 313 1318
<< polysilicon >>
rect -100 1327 100 1340
rect -100 1281 -87 1327
rect 87 1281 100 1327
rect -100 1248 100 1281
rect -100 765 100 798
rect -100 719 -87 765
rect 87 719 100 765
rect -100 706 100 719
rect -100 645 100 658
rect -100 599 -87 645
rect 87 599 100 645
rect -100 566 100 599
rect -100 83 100 116
rect -100 37 -87 83
rect 87 37 100 83
rect -100 24 100 37
rect -100 -37 100 -24
rect -100 -83 -87 -37
rect 87 -83 100 -37
rect -100 -116 100 -83
rect -100 -599 100 -566
rect -100 -645 -87 -599
rect 87 -645 100 -599
rect -100 -658 100 -645
rect -100 -719 100 -706
rect -100 -765 -87 -719
rect 87 -765 100 -719
rect -100 -798 100 -765
rect -100 -1281 100 -1248
rect -100 -1327 -87 -1281
rect 87 -1327 100 -1281
rect -100 -1340 100 -1327
<< polycontact >>
rect -87 1281 87 1327
rect -87 719 87 765
rect -87 599 87 645
rect -87 37 87 83
rect -87 -83 87 -37
rect -87 -645 87 -599
rect -87 -765 87 -719
rect -87 -1327 87 -1281
<< metal1 >>
rect -313 1375 313 1421
rect -313 1318 -267 1375
rect -98 1281 -87 1327
rect 87 1281 98 1327
rect 267 1318 313 1375
rect -175 1235 -129 1246
rect -175 800 -129 811
rect 129 1235 175 1246
rect 129 800 175 811
rect -98 719 -87 765
rect 87 719 98 765
rect -98 599 -87 645
rect 87 599 98 645
rect -175 553 -129 564
rect -175 118 -129 129
rect 129 553 175 564
rect 129 118 175 129
rect -98 37 -87 83
rect 87 37 98 83
rect -98 -83 -87 -37
rect 87 -83 98 -37
rect -175 -129 -129 -118
rect -175 -564 -129 -553
rect 129 -129 175 -118
rect 129 -564 175 -553
rect -98 -645 -87 -599
rect 87 -645 98 -599
rect -98 -765 -87 -719
rect 87 -765 98 -719
rect -175 -811 -129 -800
rect -175 -1246 -129 -1235
rect 129 -811 175 -800
rect 129 -1246 175 -1235
rect -313 -1375 -267 -1318
rect -98 -1327 -87 -1281
rect 87 -1327 98 -1281
rect 267 -1375 313 -1318
rect -313 -1421 313 -1375
<< properties >>
string FIXED_BBOX -290 -1398 290 1398
string gencell nfet_03v3
string library gf180mcu
string parameters w 2.25 l 1.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
