* Extracted by KLayout with GF180MCU LVS runset on : 05/09/2025 10:21

.SUBCKT dff_2ph_clk VSS|VSSD D D|Q Q CLK_PH2|E CLK_PH1|E VDD|VDDD gf180mcu_gnd
M$1 VDD|VDDD CLK_PH1|E \$2 VDD|VDDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P
+ AD=0.476P PS=3.64U PD=2.18U
M$2 \$3 \$2 VDD|VDDD VDD|VDDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$3 VDD|VDDD CLK_PH2|E \$8 VDD|VDDD pfet_05v0 L=0.5U W=1.38U AS=0.6072P
+ AD=0.476P PS=3.64U PD=2.18U
M$4 \$9 \$8 VDD|VDDD VDD|VDDD pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$5 \$29 D VDD|VDDD VDD|VDDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$6 \$5 \$2 \$29 VDD|VDDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$7 \$5 \$3 \$30 VDD|VDDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$8 VDD|VDDD \$6 \$30 VDD|VDDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$9 \$6 \$5 VDD|VDDD VDD|VDDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$10 \$36 D|Q VDD|VDDD VDD|VDDD pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$11 \$10 \$8 \$36 VDD|VDDD pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$12 \$10 \$9 \$37 VDD|VDDD pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$13 VDD|VDDD \$11 \$37 VDD|VDDD pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$14 \$11 \$10 VDD|VDDD VDD|VDDD pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$15 VDD|VDDD \$5 D|Q VDD|VDDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$16 VDD|VDDD \$10 Q VDD|VDDD pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$17 \$19 D VSS|VSSD gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$18 \$5 \$3 \$19 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$19 \$18 \$2 \$5 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$20 VSS|VSSD \$6 \$18 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.263P
+ AD=0.2054P PS=1.49U PD=1.31U
M$21 \$6 \$5 VSS|VSSD gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.2054P
+ AD=0.3476P PS=1.31U PD=2.46U
M$22 \$26 D|Q VSS|VSSD gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P
+ PS=2.28U PD=0.94U
M$23 \$10 \$9 \$26 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P
+ PS=0.94U PD=1.22U
M$24 \$23 \$8 \$10 gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P
+ PS=1.22U PD=1.49U
M$25 VSS|VSSD \$11 \$23 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.263P
+ AD=0.2054P PS=1.49U PD=1.31U
M$26 \$11 \$10 VSS|VSSD gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.2054P
+ AD=0.3476P PS=1.31U PD=2.46U
M$27 VSS|VSSD CLK_PH1|E \$2 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.3476P
+ AD=0.263P PS=2.46U PD=1.49U
M$28 \$3 \$2 VSS|VSSD gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$29 VSS|VSSD CLK_PH2|E \$8 gf180mcu_gnd nfet_05v0 L=0.6U W=0.79U AS=0.3476P
+ AD=0.263P PS=2.46U PD=1.49U
M$30 \$9 \$8 VSS|VSSD gf180mcu_gnd nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P
+ PS=1.49U PD=2.28U
M$31 VSS|VSSD \$5 D|Q gf180mcu_gnd nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
M$32 VSS|VSSD \$10 Q gf180mcu_gnd nfet_05v0 L=0.6U W=1.32U AS=0.5808P
+ AD=0.5808P PS=3.52U PD=3.52U
.ENDS dff_2ph_clk
