magic
tech gf180mcuD
magscale 1 10
timestamp 1757672677
<< error_s >>
rect 315 -1058 317 -798
<< metal1 >>
rect -1224 1370 2180 1570
rect -1224 274 -1124 1370
rect -920 388 1876 400
rect -920 336 -126 388
rect -74 336 1876 388
rect -920 324 1876 336
rect 2080 274 2180 1370
rect -1224 174 2180 274
rect -1171 -110 -991 174
rect 423 -110 603 174
rect -1171 -290 603 -110
rect 704 -24 2172 76
rect -661 -726 -613 -702
rect -625 -778 -613 -726
rect -661 -802 -613 -778
rect -386 -726 -245 -702
rect -386 -778 -374 -726
rect -386 -802 -245 -778
rect -68 -802 203 -702
rect 704 -1118 804 -24
rect 1000 -1004 1876 -992
rect 1000 -1056 1012 -1004
rect 1064 -1056 1172 -1004
rect 1224 -1056 1332 -1004
rect 1384 -1056 1492 -1004
rect 1544 -1056 1652 -1004
rect 1704 -1056 1812 -1004
rect 1864 -1056 1876 -1004
rect 1000 -1068 1876 -1056
rect 2072 -1118 2172 -24
rect -1224 -1318 2180 -1118
<< via1 >>
rect -1020 574 -968 1146
rect -828 574 -776 1146
rect -668 574 -616 1146
rect -508 574 -456 1146
rect -348 574 -296 1146
rect -188 574 -136 1146
rect -28 574 24 1146
rect 132 574 184 1146
rect 292 574 344 1146
rect 452 574 504 1146
rect 612 574 664 1146
rect 772 574 824 1146
rect 932 574 984 1146
rect 1092 574 1144 1146
rect 1252 574 1304 1146
rect 1412 574 1464 1146
rect 1572 574 1624 1146
rect 1732 574 1784 1146
rect 1924 574 1976 1146
rect -126 336 -74 388
rect -1036 -834 -984 -678
rect -805 -722 -753 -566
rect -677 -778 -625 -726
rect -374 -778 -218 -726
rect -126 -1058 -74 -798
rect 315 -1058 367 -798
rect 904 -820 956 -248
rect 1092 -820 1144 -248
rect 1252 -820 1304 -248
rect 1412 -820 1464 -248
rect 1572 -820 1624 -248
rect 1732 -820 1784 -248
rect 1920 -820 1972 -248
rect 1012 -1056 1064 -1004
rect 1172 -1056 1224 -1004
rect 1332 -1056 1384 -1004
rect 1492 -1056 1544 -1004
rect 1652 -1056 1704 -1004
rect 1812 -1056 1864 -1004
<< metal2 >>
rect -1032 1146 -924 1284
rect -1032 976 -1020 1146
rect -968 976 -924 1146
rect -1032 920 -1022 976
rect -966 920 -924 976
rect -1032 852 -1020 920
rect -968 852 -924 920
rect -1032 796 -1022 852
rect -966 796 -924 852
rect -1032 574 -1020 796
rect -968 574 -924 796
rect -1032 516 -924 574
rect -840 1274 -764 1284
rect -840 1218 -829 1274
rect -773 1218 -764 1274
rect -840 1150 -764 1218
rect -840 1094 -829 1150
rect -773 1094 -764 1150
rect -840 574 -828 1094
rect -776 574 -764 1094
rect -840 516 -764 574
rect -680 1146 -604 1284
rect -680 976 -668 1146
rect -616 976 -604 1146
rect -680 920 -670 976
rect -614 920 -604 976
rect -680 852 -668 920
rect -616 852 -604 920
rect -680 796 -670 852
rect -614 796 -604 852
rect -680 574 -668 796
rect -616 574 -604 796
rect -680 516 -604 574
rect -520 1274 -444 1284
rect -520 1218 -510 1274
rect -454 1218 -444 1274
rect -520 1150 -444 1218
rect -520 1094 -510 1150
rect -454 1094 -444 1150
rect -520 574 -508 1094
rect -456 574 -444 1094
rect -520 516 -444 574
rect -360 1146 -284 1284
rect -360 976 -348 1146
rect -296 976 -284 1146
rect -360 920 -350 976
rect -294 920 -284 976
rect -360 852 -348 920
rect -296 852 -284 920
rect -360 796 -350 852
rect -294 796 -284 852
rect -360 574 -348 796
rect -296 574 -284 796
rect -360 516 -284 574
rect -200 1274 -124 1284
rect -200 1218 -190 1274
rect -134 1218 -124 1274
rect -200 1150 -124 1218
rect -200 1094 -190 1150
rect -134 1094 -124 1150
rect -200 574 -188 1094
rect -136 574 -124 1094
rect -200 516 -124 574
rect -40 1146 36 1284
rect -40 976 -28 1146
rect 24 976 36 1146
rect -40 920 -30 976
rect 26 920 36 976
rect -40 852 -28 920
rect 24 852 36 920
rect -40 796 -30 852
rect 26 796 36 852
rect -40 574 -28 796
rect 24 574 36 796
rect -40 516 36 574
rect 120 1274 196 1284
rect 120 1218 131 1274
rect 187 1218 196 1274
rect 120 1150 196 1218
rect 120 1094 131 1150
rect 187 1094 196 1150
rect 120 574 132 1094
rect 184 574 196 1094
rect 120 516 196 574
rect 280 1146 356 1284
rect 280 976 292 1146
rect 344 976 356 1146
rect 280 920 290 976
rect 346 920 356 976
rect 280 852 292 920
rect 344 852 356 920
rect 280 796 290 852
rect 346 796 356 852
rect 280 574 292 796
rect 344 574 356 796
rect 280 516 356 574
rect 440 1274 516 1284
rect 440 1218 450 1274
rect 506 1218 516 1274
rect 440 1150 516 1218
rect 440 1094 450 1150
rect 506 1094 516 1150
rect 440 574 452 1094
rect 504 574 516 1094
rect 440 516 516 574
rect 600 1146 676 1284
rect 600 976 612 1146
rect 664 976 676 1146
rect 600 920 610 976
rect 666 920 676 976
rect 600 852 612 920
rect 664 852 676 920
rect 600 796 610 852
rect 666 796 676 852
rect 600 574 612 796
rect 664 574 676 796
rect 600 516 676 574
rect 760 1274 836 1284
rect 760 1218 770 1274
rect 826 1218 836 1274
rect 760 1150 836 1218
rect 760 1094 770 1150
rect 826 1094 836 1150
rect 760 574 772 1094
rect 824 574 836 1094
rect 760 516 836 574
rect 920 1146 996 1284
rect 920 976 932 1146
rect 984 976 996 1146
rect 920 920 930 976
rect 986 920 996 976
rect 920 852 932 920
rect 984 852 996 920
rect 920 796 930 852
rect 986 796 996 852
rect 920 574 932 796
rect 984 574 996 796
rect -150 388 -50 400
rect -150 336 -126 388
rect -74 336 -50 388
rect -845 -366 -745 -356
rect -845 -422 -823 -366
rect -767 -422 -745 -366
rect -1060 -522 -960 -512
rect -1060 -578 -1038 -522
rect -982 -578 -960 -522
rect -1060 -678 -960 -578
rect -1060 -834 -1036 -678
rect -984 -834 -960 -678
rect -845 -566 -745 -422
rect -845 -722 -805 -566
rect -753 -722 -745 -566
rect -845 -734 -745 -722
rect -689 -726 -206 -702
rect -689 -778 -677 -726
rect -625 -778 -374 -726
rect -218 -778 -206 -726
rect -689 -802 -206 -778
rect -150 -798 -50 336
rect 920 -190 996 574
rect 892 -248 996 -190
rect -1060 -846 -960 -834
rect -150 -1058 -126 -798
rect -74 -1058 -50 -798
rect -150 -1072 -50 -1058
rect 315 -798 415 -786
rect 367 -980 415 -798
rect 892 -820 904 -248
rect 956 -820 996 -248
rect 892 -878 996 -820
rect 1080 1274 1156 1284
rect 1080 1218 1091 1274
rect 1147 1218 1156 1274
rect 1080 1150 1156 1218
rect 1080 1094 1091 1150
rect 1147 1094 1156 1150
rect 1080 574 1092 1094
rect 1144 574 1156 1094
rect 1080 -248 1156 574
rect 1080 -820 1092 -248
rect 1144 -820 1156 -248
rect 1080 -878 1156 -820
rect 1240 1146 1316 1284
rect 1240 976 1252 1146
rect 1304 976 1316 1146
rect 1240 920 1250 976
rect 1306 920 1316 976
rect 1240 852 1252 920
rect 1304 852 1316 920
rect 1240 796 1250 852
rect 1306 796 1316 852
rect 1240 574 1252 796
rect 1304 574 1316 796
rect 1240 -248 1316 574
rect 1240 -820 1252 -248
rect 1304 -820 1316 -248
rect 1240 -878 1316 -820
rect 1400 1274 1476 1284
rect 1400 1218 1410 1274
rect 1466 1218 1476 1274
rect 1400 1150 1476 1218
rect 1400 1094 1410 1150
rect 1466 1094 1476 1150
rect 1400 574 1412 1094
rect 1464 574 1476 1094
rect 1400 -248 1476 574
rect 1400 -820 1412 -248
rect 1464 -820 1476 -248
rect 1400 -878 1476 -820
rect 1560 1146 1636 1284
rect 1560 976 1572 1146
rect 1624 976 1636 1146
rect 1560 920 1570 976
rect 1626 920 1636 976
rect 1560 852 1572 920
rect 1624 852 1636 920
rect 1560 796 1570 852
rect 1626 796 1636 852
rect 1560 574 1572 796
rect 1624 574 1636 796
rect 1560 -248 1636 574
rect 1560 -820 1572 -248
rect 1624 -820 1636 -248
rect 1560 -878 1636 -820
rect 1720 1274 1796 1284
rect 1720 1218 1730 1274
rect 1786 1218 1796 1274
rect 1720 1150 1796 1218
rect 1720 1094 1730 1150
rect 1786 1094 1796 1150
rect 1720 574 1732 1094
rect 1784 574 1796 1094
rect 1720 -248 1796 574
rect 1720 -820 1732 -248
rect 1784 -820 1796 -248
rect 1720 -878 1796 -820
rect 1880 1146 1988 1284
rect 1880 976 1924 1146
rect 1976 976 1988 1146
rect 1880 920 1922 976
rect 1978 920 1988 976
rect 1880 852 1924 920
rect 1976 852 1988 920
rect 1880 796 1922 852
rect 1978 796 1988 852
rect 1880 574 1924 796
rect 1976 574 1988 796
rect 1880 516 1988 574
rect 1880 -190 1956 516
rect 1880 -248 1984 -190
rect 1880 -820 1920 -248
rect 1972 -820 1984 -248
rect 1880 -878 1984 -820
rect 367 -1004 1876 -980
rect 367 -1056 1012 -1004
rect 1064 -1056 1172 -1004
rect 1224 -1056 1332 -1004
rect 1384 -1056 1492 -1004
rect 1544 -1056 1652 -1004
rect 1704 -1056 1812 -1004
rect 1864 -1056 1876 -1004
rect 367 -1058 1876 -1056
rect 315 -1080 1876 -1058
<< via2 >>
rect -1022 920 -1020 976
rect -1020 920 -968 976
rect -968 920 -966 976
rect -1022 796 -1020 852
rect -1020 796 -968 852
rect -968 796 -966 852
rect -829 1218 -773 1274
rect -829 1146 -773 1150
rect -829 1094 -828 1146
rect -828 1094 -776 1146
rect -776 1094 -773 1146
rect -670 920 -668 976
rect -668 920 -616 976
rect -616 920 -614 976
rect -670 796 -668 852
rect -668 796 -616 852
rect -616 796 -614 852
rect -510 1218 -454 1274
rect -510 1146 -454 1150
rect -510 1094 -508 1146
rect -508 1094 -456 1146
rect -456 1094 -454 1146
rect -350 920 -348 976
rect -348 920 -296 976
rect -296 920 -294 976
rect -350 796 -348 852
rect -348 796 -296 852
rect -296 796 -294 852
rect -190 1218 -134 1274
rect -190 1146 -134 1150
rect -190 1094 -188 1146
rect -188 1094 -136 1146
rect -136 1094 -134 1146
rect -30 920 -28 976
rect -28 920 24 976
rect 24 920 26 976
rect -30 796 -28 852
rect -28 796 24 852
rect 24 796 26 852
rect 131 1218 187 1274
rect 131 1146 187 1150
rect 131 1094 132 1146
rect 132 1094 184 1146
rect 184 1094 187 1146
rect 290 920 292 976
rect 292 920 344 976
rect 344 920 346 976
rect 290 796 292 852
rect 292 796 344 852
rect 344 796 346 852
rect 450 1218 506 1274
rect 450 1146 506 1150
rect 450 1094 452 1146
rect 452 1094 504 1146
rect 504 1094 506 1146
rect 610 920 612 976
rect 612 920 664 976
rect 664 920 666 976
rect 610 796 612 852
rect 612 796 664 852
rect 664 796 666 852
rect 770 1218 826 1274
rect 770 1146 826 1150
rect 770 1094 772 1146
rect 772 1094 824 1146
rect 824 1094 826 1146
rect 930 920 932 976
rect 932 920 984 976
rect 984 920 986 976
rect 930 796 932 852
rect 932 796 984 852
rect 984 796 986 852
rect -823 -422 -767 -366
rect -1038 -578 -982 -522
rect 1091 1218 1147 1274
rect 1091 1146 1147 1150
rect 1091 1094 1092 1146
rect 1092 1094 1144 1146
rect 1144 1094 1147 1146
rect 1250 920 1252 976
rect 1252 920 1304 976
rect 1304 920 1306 976
rect 1250 796 1252 852
rect 1252 796 1304 852
rect 1304 796 1306 852
rect 1410 1218 1466 1274
rect 1410 1146 1466 1150
rect 1410 1094 1412 1146
rect 1412 1094 1464 1146
rect 1464 1094 1466 1146
rect 1570 920 1572 976
rect 1572 920 1624 976
rect 1624 920 1626 976
rect 1570 796 1572 852
rect 1572 796 1624 852
rect 1624 796 1626 852
rect 1730 1218 1786 1274
rect 1730 1146 1786 1150
rect 1730 1094 1732 1146
rect 1732 1094 1784 1146
rect 1784 1094 1786 1146
rect 1922 920 1924 976
rect 1924 920 1976 976
rect 1976 920 1978 976
rect 1922 796 1924 852
rect 1924 796 1976 852
rect 1976 796 1978 852
<< metal3 >>
rect -1224 1274 2080 1284
rect -1224 1218 -829 1274
rect -773 1218 -510 1274
rect -454 1218 -190 1274
rect -134 1218 131 1274
rect 187 1218 450 1274
rect 506 1218 770 1274
rect 826 1218 1091 1274
rect 1147 1218 1410 1274
rect 1466 1218 1730 1274
rect 1786 1218 2080 1274
rect -1224 1150 2080 1218
rect -1224 1094 -829 1150
rect -773 1094 -510 1150
rect -454 1094 -190 1150
rect -134 1094 131 1150
rect 187 1094 450 1150
rect 506 1094 770 1150
rect 826 1094 1091 1150
rect 1147 1094 1410 1150
rect 1466 1094 1730 1150
rect 1786 1094 2080 1150
rect -1224 1084 2080 1094
rect -1224 976 2080 986
rect -1224 920 -1022 976
rect -966 920 -670 976
rect -614 920 -350 976
rect -294 920 -30 976
rect 26 920 290 976
rect 346 920 610 976
rect 666 920 930 976
rect 986 920 1250 976
rect 1306 920 1570 976
rect 1626 920 1922 976
rect 1978 920 2080 976
rect -1224 852 2080 920
rect -1224 796 -1022 852
rect -966 796 -670 852
rect -614 796 -350 852
rect -294 796 -30 852
rect 26 796 290 852
rect 346 796 610 852
rect 666 796 930 852
rect 986 796 1250 852
rect 1306 796 1570 852
rect 1626 796 1922 852
rect 1978 796 2080 852
rect -1224 786 2080 796
rect -1171 -366 -745 -344
rect -1171 -422 -823 -366
rect -767 -422 -745 -366
rect -1171 -444 -745 -422
rect -1171 -522 2180 -500
rect -1171 -578 -1038 -522
rect -982 -578 2180 -522
rect -1171 -600 2180 -578
use gf180mcu_fd_sc_mcu9t5v0__filltie  gf180mcu_fd_sc_mcu9t5v0__filltie_0
timestamp 1757672677
transform 1 0 -611 0 1 -1208
box -86 -90 310 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  gf180mcu_fd_sc_mcu9t5v0__inv_1_0
timestamp 1757672677
transform 1 0 -387 0 1 -1208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__inv_1  gf180mcu_fd_sc_mcu9t5v0__inv_1_1
timestamp 1757672677
transform 1 0 61 0 1 -1208
box -86 -90 534 1098
use gf180mcu_fd_sc_mcu9t5v0__nand2_1  gf180mcu_fd_sc_mcu9t5v0__nand2_1_0
timestamp 1757672677
transform 1 0 -1171 0 1 -1208
box -86 -90 646 1098
use nfet  nfet_0
timestamp 1757672677
transform 1 0 972 0 1 -934
box -268 -284 1200 1010
use pfet  pfet_0
timestamp 1757672677
transform 1 0 -948 0 1 460
box -352 -362 3204 1086
<< labels >>
flabel metal1 s -1168 1567 -1168 1567 4 FreeSans 73 0 0 0 VDDD
port 1 nsew
flabel metal1 s 608 1567 608 1567 4 FreeSans 73 0 0 0 VDDD
port 1 nsew
flabel metal1 s -1168 -1295 -1168 -1295 2 FreeSans 73 0 0 0 VSSD
port 2 nsew
flabel metal1 s 606 -1315 606 -1315 2 FreeSans 73 0 0 0 VSSD
port 2 nsew
flabel metal3 s -1168 1184 -1168 1184 2 FreeSans 89 0 0 0 T1
port 3 nsew
flabel metal3 s -1168 886 -1168 886 2 FreeSans 89 0 0 0 T2
port 4 nsew
flabel metal3 s -1168 -394 -1168 -394 2 FreeSans 89 0 0 0 CON
port 5 nsew
flabel metal3 s -1168 -550 -1168 -550 2 FreeSans 89 0 0 0 EN
port 6 nsew
<< properties >>
string path 10.400 5.920 -6.120 5.920 
<< end >>
