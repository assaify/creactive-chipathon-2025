magic
tech gf180mcuD
magscale 1 10
timestamp 1755276408
<< pwell >>
rect -350 -2458 350 2458
<< nmos >>
rect -100 1298 100 2248
rect -100 116 100 1066
rect -100 -1066 100 -116
rect -100 -2248 100 -1298
<< ndiff >>
rect -188 2235 -100 2248
rect -188 1311 -175 2235
rect -129 1311 -100 2235
rect -188 1298 -100 1311
rect 100 2235 188 2248
rect 100 1311 129 2235
rect 175 1311 188 2235
rect 100 1298 188 1311
rect -188 1053 -100 1066
rect -188 129 -175 1053
rect -129 129 -100 1053
rect -188 116 -100 129
rect 100 1053 188 1066
rect 100 129 129 1053
rect 175 129 188 1053
rect 100 116 188 129
rect -188 -129 -100 -116
rect -188 -1053 -175 -129
rect -129 -1053 -100 -129
rect -188 -1066 -100 -1053
rect 100 -129 188 -116
rect 100 -1053 129 -129
rect 175 -1053 188 -129
rect 100 -1066 188 -1053
rect -188 -1311 -100 -1298
rect -188 -2235 -175 -1311
rect -129 -2235 -100 -1311
rect -188 -2248 -100 -2235
rect 100 -1311 188 -1298
rect 100 -2235 129 -1311
rect 175 -2235 188 -1311
rect 100 -2248 188 -2235
<< ndiffc >>
rect -175 1311 -129 2235
rect 129 1311 175 2235
rect -175 129 -129 1053
rect 129 129 175 1053
rect -175 -1053 -129 -129
rect 129 -1053 175 -129
rect -175 -2235 -129 -1311
rect 129 -2235 175 -1311
<< psubdiff >>
rect -326 2362 326 2434
rect -326 2318 -254 2362
rect -326 -2318 -313 2318
rect -267 -2318 -254 2318
rect 254 2318 326 2362
rect -326 -2362 -254 -2318
rect 254 -2318 267 2318
rect 313 -2318 326 2318
rect 254 -2362 326 -2318
rect -326 -2434 326 -2362
<< psubdiffcont >>
rect -313 -2318 -267 2318
rect 267 -2318 313 2318
<< polysilicon >>
rect -100 2327 100 2340
rect -100 2281 -87 2327
rect 87 2281 100 2327
rect -100 2248 100 2281
rect -100 1265 100 1298
rect -100 1219 -87 1265
rect 87 1219 100 1265
rect -100 1206 100 1219
rect -100 1145 100 1158
rect -100 1099 -87 1145
rect 87 1099 100 1145
rect -100 1066 100 1099
rect -100 83 100 116
rect -100 37 -87 83
rect 87 37 100 83
rect -100 24 100 37
rect -100 -37 100 -24
rect -100 -83 -87 -37
rect 87 -83 100 -37
rect -100 -116 100 -83
rect -100 -1099 100 -1066
rect -100 -1145 -87 -1099
rect 87 -1145 100 -1099
rect -100 -1158 100 -1145
rect -100 -1219 100 -1206
rect -100 -1265 -87 -1219
rect 87 -1265 100 -1219
rect -100 -1298 100 -1265
rect -100 -2281 100 -2248
rect -100 -2327 -87 -2281
rect 87 -2327 100 -2281
rect -100 -2340 100 -2327
<< polycontact >>
rect -87 2281 87 2327
rect -87 1219 87 1265
rect -87 1099 87 1145
rect -87 37 87 83
rect -87 -83 87 -37
rect -87 -1145 87 -1099
rect -87 -1265 87 -1219
rect -87 -2327 87 -2281
<< metal1 >>
rect -313 2375 313 2421
rect -313 2318 -267 2375
rect -98 2281 -87 2327
rect 87 2281 98 2327
rect 267 2318 313 2375
rect -175 2235 -129 2246
rect -175 1300 -129 1311
rect 129 2235 175 2246
rect 129 1300 175 1311
rect -98 1219 -87 1265
rect 87 1219 98 1265
rect -98 1099 -87 1145
rect 87 1099 98 1145
rect -175 1053 -129 1064
rect -175 118 -129 129
rect 129 1053 175 1064
rect 129 118 175 129
rect -98 37 -87 83
rect 87 37 98 83
rect -98 -83 -87 -37
rect 87 -83 98 -37
rect -175 -129 -129 -118
rect -175 -1064 -129 -1053
rect 129 -129 175 -118
rect 129 -1064 175 -1053
rect -98 -1145 -87 -1099
rect 87 -1145 98 -1099
rect -98 -1265 -87 -1219
rect 87 -1265 98 -1219
rect -175 -1311 -129 -1300
rect -175 -2246 -129 -2235
rect 129 -1311 175 -1300
rect 129 -2246 175 -2235
rect -313 -2375 -267 -2318
rect -98 -2327 -87 -2281
rect 87 -2327 98 -2281
rect 267 -2375 313 -2318
rect -313 -2421 313 -2375
<< properties >>
string FIXED_BBOX -290 -2398 290 2398
string gencell nfet_03v3
string library gf180mcu
string parameters w 4.75 l 1.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
