magic
tech gf180mcuD
magscale 1 10
timestamp 1755277289
<< pwell >>
rect -1596 -1695 1596 1695
<< psubdiff >>
rect -1572 1599 1572 1671
rect -1572 1555 -1500 1599
rect -1572 -1555 -1559 1555
rect -1513 -1555 -1500 1555
rect 1500 1555 1572 1599
rect -1572 -1599 -1500 -1555
rect 1500 -1555 1513 1555
rect 1559 -1555 1572 1555
rect 1500 -1599 1572 -1555
rect -1572 -1671 1572 -1599
<< psubdiffcont >>
rect -1559 -1555 -1513 1555
rect 1513 -1555 1559 1555
<< polysilicon >>
rect -1360 1446 -1160 1459
rect -1360 1400 -1347 1446
rect -1173 1400 -1160 1446
rect -1360 1337 -1160 1400
rect -1360 -1400 -1160 -1337
rect -1360 -1446 -1347 -1400
rect -1173 -1446 -1160 -1400
rect -1360 -1459 -1160 -1446
rect -1080 1446 -880 1459
rect -1080 1400 -1067 1446
rect -893 1400 -880 1446
rect -1080 1337 -880 1400
rect -1080 -1400 -880 -1337
rect -1080 -1446 -1067 -1400
rect -893 -1446 -880 -1400
rect -1080 -1459 -880 -1446
rect -800 1446 -600 1459
rect -800 1400 -787 1446
rect -613 1400 -600 1446
rect -800 1337 -600 1400
rect -800 -1400 -600 -1337
rect -800 -1446 -787 -1400
rect -613 -1446 -600 -1400
rect -800 -1459 -600 -1446
rect -520 1446 -320 1459
rect -520 1400 -507 1446
rect -333 1400 -320 1446
rect -520 1337 -320 1400
rect -520 -1400 -320 -1337
rect -520 -1446 -507 -1400
rect -333 -1446 -320 -1400
rect -520 -1459 -320 -1446
rect -240 1446 -40 1459
rect -240 1400 -227 1446
rect -53 1400 -40 1446
rect -240 1337 -40 1400
rect -240 -1400 -40 -1337
rect -240 -1446 -227 -1400
rect -53 -1446 -40 -1400
rect -240 -1459 -40 -1446
rect 40 1446 240 1459
rect 40 1400 53 1446
rect 227 1400 240 1446
rect 40 1337 240 1400
rect 40 -1400 240 -1337
rect 40 -1446 53 -1400
rect 227 -1446 240 -1400
rect 40 -1459 240 -1446
rect 320 1446 520 1459
rect 320 1400 333 1446
rect 507 1400 520 1446
rect 320 1337 520 1400
rect 320 -1400 520 -1337
rect 320 -1446 333 -1400
rect 507 -1446 520 -1400
rect 320 -1459 520 -1446
rect 600 1446 800 1459
rect 600 1400 613 1446
rect 787 1400 800 1446
rect 600 1337 800 1400
rect 600 -1400 800 -1337
rect 600 -1446 613 -1400
rect 787 -1446 800 -1400
rect 600 -1459 800 -1446
rect 880 1446 1080 1459
rect 880 1400 893 1446
rect 1067 1400 1080 1446
rect 880 1337 1080 1400
rect 880 -1400 1080 -1337
rect 880 -1446 893 -1400
rect 1067 -1446 1080 -1400
rect 880 -1459 1080 -1446
rect 1160 1446 1360 1459
rect 1160 1400 1173 1446
rect 1347 1400 1360 1446
rect 1160 1337 1360 1400
rect 1160 -1400 1360 -1337
rect 1160 -1446 1173 -1400
rect 1347 -1446 1360 -1400
rect 1160 -1459 1360 -1446
<< polycontact >>
rect -1347 1400 -1173 1446
rect -1347 -1446 -1173 -1400
rect -1067 1400 -893 1446
rect -1067 -1446 -893 -1400
rect -787 1400 -613 1446
rect -787 -1446 -613 -1400
rect -507 1400 -333 1446
rect -507 -1446 -333 -1400
rect -227 1400 -53 1446
rect -227 -1446 -53 -1400
rect 53 1400 227 1446
rect 53 -1446 227 -1400
rect 333 1400 507 1446
rect 333 -1446 507 -1400
rect 613 1400 787 1446
rect 613 -1446 787 -1400
rect 893 1400 1067 1446
rect 893 -1446 1067 -1400
rect 1173 1400 1347 1446
rect 1173 -1446 1347 -1400
<< nhighres >>
rect -1360 -1337 -1160 1337
rect -1080 -1337 -880 1337
rect -800 -1337 -600 1337
rect -520 -1337 -320 1337
rect -240 -1337 -40 1337
rect 40 -1337 240 1337
rect 320 -1337 520 1337
rect 600 -1337 800 1337
rect 880 -1337 1080 1337
rect 1160 -1337 1360 1337
<< metal1 >>
rect -1559 1612 1559 1658
rect -1559 1555 -1513 1612
rect 1513 1555 1559 1612
rect -1358 1400 -1347 1446
rect -1173 1400 -1162 1446
rect -1078 1400 -1067 1446
rect -893 1400 -882 1446
rect -798 1400 -787 1446
rect -613 1400 -602 1446
rect -518 1400 -507 1446
rect -333 1400 -322 1446
rect -238 1400 -227 1446
rect -53 1400 -42 1446
rect 42 1400 53 1446
rect 227 1400 238 1446
rect 322 1400 333 1446
rect 507 1400 518 1446
rect 602 1400 613 1446
rect 787 1400 798 1446
rect 882 1400 893 1446
rect 1067 1400 1078 1446
rect 1162 1400 1173 1446
rect 1347 1400 1358 1446
rect -1358 -1446 -1347 -1400
rect -1173 -1446 -1162 -1400
rect -1078 -1446 -1067 -1400
rect -893 -1446 -882 -1400
rect -798 -1446 -787 -1400
rect -613 -1446 -602 -1400
rect -518 -1446 -507 -1400
rect -333 -1446 -322 -1400
rect -238 -1446 -227 -1400
rect -53 -1446 -42 -1400
rect 42 -1446 53 -1400
rect 227 -1446 238 -1400
rect 322 -1446 333 -1400
rect 507 -1446 518 -1400
rect 602 -1446 613 -1400
rect 787 -1446 798 -1400
rect 882 -1446 893 -1400
rect 1067 -1446 1078 -1400
rect 1162 -1446 1173 -1400
rect 1347 -1446 1358 -1400
rect -1559 -1612 -1513 -1555
rect 1513 -1612 1559 -1555
rect -1559 -1658 1559 -1612
<< properties >>
string FIXED_BBOX -1536 -1635 1536 1635
string gencell ppolyf_u_1k
string library gf180mcu
string parameters w 1.0 l 13.37 m 1 nx 10 wmin 1.000 lmin 1.000 class resistor rho 1000 val 13.37k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
