* Extracted by KLayout with GF180MCU LVS runset on : 04/09/2025 15:13

.SUBCKT tail_current VSS I2A I1C I1B IBIAS I2B I2C I1A
M$1 VSS VSS VSS VSS nfet_03v3 L=0.8U W=105U AS=45.15P AD=45.15P PS=144.08U
+ PD=144.08U
M$2 I2A IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$12 I1C IBIAS VSS VSS nfet_03v3 L=0.8U W=7.5U AS=3P AD=3P PS=9.1U PD=9.1U
M$13 I1C I1C I1C VSS nfet_03v3 L=0.8U W=7.5U AS=3.7875P AD=3.7875P PS=13.27U
+ PD=13.27U
M$14 I1B I1B I1B VSS nfet_03v3 L=0.8U W=7.5U AS=3.7875P AD=3.7875P PS=13.27U
+ PD=13.27U
M$15 VSS IBIAS I1B VSS nfet_03v3 L=0.8U W=7.5U AS=3P AD=3P PS=9.1U PD=9.1U
M$28 I2B IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$30 I2C IBIAS VSS VSS nfet_03v3 L=0.8U W=75U AS=30P AD=30P PS=91U PD=91U
M$38 I1A IBIAS VSS VSS nfet_03v3 L=0.8U W=7.5U AS=3P AD=3P PS=9.1U PD=9.1U
M$39 I1A I1A I1A VSS nfet_03v3 L=0.8U W=7.5U AS=3.7875P AD=3.7875P PS=13.27U
+ PD=13.27U
M$40 IBIAS IBIAS IBIAS VSS nfet_03v3 L=0.8U W=7.5U AS=3.7875P AD=3.7875P
+ PS=13.27U PD=13.27U
M$41 VSS IBIAS IBIAS VSS nfet_03v3 L=0.8U W=7.5U AS=3P AD=3P PS=9.1U PD=9.1U
.ENDS tail_current
