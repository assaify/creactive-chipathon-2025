magic
tech gf180mcuD
magscale 1 10
timestamp 1755277289
<< pwell >>
rect -3238 -435 3238 435
<< nmos >>
rect -2988 -225 -2788 225
rect -2684 -225 -2484 225
rect -2380 -225 -2180 225
rect -2076 -225 -1876 225
rect -1772 -225 -1572 225
rect -1468 -225 -1268 225
rect -1164 -225 -964 225
rect -860 -225 -660 225
rect -556 -225 -356 225
rect -252 -225 -52 225
rect 52 -225 252 225
rect 356 -225 556 225
rect 660 -225 860 225
rect 964 -225 1164 225
rect 1268 -225 1468 225
rect 1572 -225 1772 225
rect 1876 -225 2076 225
rect 2180 -225 2380 225
rect 2484 -225 2684 225
rect 2788 -225 2988 225
<< ndiff >>
rect -3076 212 -2988 225
rect -3076 -212 -3063 212
rect -3017 -212 -2988 212
rect -3076 -225 -2988 -212
rect -2788 212 -2684 225
rect -2788 -212 -2759 212
rect -2713 -212 -2684 212
rect -2788 -225 -2684 -212
rect -2484 212 -2380 225
rect -2484 -212 -2455 212
rect -2409 -212 -2380 212
rect -2484 -225 -2380 -212
rect -2180 212 -2076 225
rect -2180 -212 -2151 212
rect -2105 -212 -2076 212
rect -2180 -225 -2076 -212
rect -1876 212 -1772 225
rect -1876 -212 -1847 212
rect -1801 -212 -1772 212
rect -1876 -225 -1772 -212
rect -1572 212 -1468 225
rect -1572 -212 -1543 212
rect -1497 -212 -1468 212
rect -1572 -225 -1468 -212
rect -1268 212 -1164 225
rect -1268 -212 -1239 212
rect -1193 -212 -1164 212
rect -1268 -225 -1164 -212
rect -964 212 -860 225
rect -964 -212 -935 212
rect -889 -212 -860 212
rect -964 -225 -860 -212
rect -660 212 -556 225
rect -660 -212 -631 212
rect -585 -212 -556 212
rect -660 -225 -556 -212
rect -356 212 -252 225
rect -356 -212 -327 212
rect -281 -212 -252 212
rect -356 -225 -252 -212
rect -52 212 52 225
rect -52 -212 -23 212
rect 23 -212 52 212
rect -52 -225 52 -212
rect 252 212 356 225
rect 252 -212 281 212
rect 327 -212 356 212
rect 252 -225 356 -212
rect 556 212 660 225
rect 556 -212 585 212
rect 631 -212 660 212
rect 556 -225 660 -212
rect 860 212 964 225
rect 860 -212 889 212
rect 935 -212 964 212
rect 860 -225 964 -212
rect 1164 212 1268 225
rect 1164 -212 1193 212
rect 1239 -212 1268 212
rect 1164 -225 1268 -212
rect 1468 212 1572 225
rect 1468 -212 1497 212
rect 1543 -212 1572 212
rect 1468 -225 1572 -212
rect 1772 212 1876 225
rect 1772 -212 1801 212
rect 1847 -212 1876 212
rect 1772 -225 1876 -212
rect 2076 212 2180 225
rect 2076 -212 2105 212
rect 2151 -212 2180 212
rect 2076 -225 2180 -212
rect 2380 212 2484 225
rect 2380 -212 2409 212
rect 2455 -212 2484 212
rect 2380 -225 2484 -212
rect 2684 212 2788 225
rect 2684 -212 2713 212
rect 2759 -212 2788 212
rect 2684 -225 2788 -212
rect 2988 212 3076 225
rect 2988 -212 3017 212
rect 3063 -212 3076 212
rect 2988 -225 3076 -212
<< ndiffc >>
rect -3063 -212 -3017 212
rect -2759 -212 -2713 212
rect -2455 -212 -2409 212
rect -2151 -212 -2105 212
rect -1847 -212 -1801 212
rect -1543 -212 -1497 212
rect -1239 -212 -1193 212
rect -935 -212 -889 212
rect -631 -212 -585 212
rect -327 -212 -281 212
rect -23 -212 23 212
rect 281 -212 327 212
rect 585 -212 631 212
rect 889 -212 935 212
rect 1193 -212 1239 212
rect 1497 -212 1543 212
rect 1801 -212 1847 212
rect 2105 -212 2151 212
rect 2409 -212 2455 212
rect 2713 -212 2759 212
rect 3017 -212 3063 212
<< psubdiff >>
rect -3214 339 3214 411
rect -3214 295 -3142 339
rect -3214 -295 -3201 295
rect -3155 -295 -3142 295
rect 3142 295 3214 339
rect -3214 -339 -3142 -295
rect 3142 -295 3155 295
rect 3201 -295 3214 295
rect 3142 -339 3214 -295
rect -3214 -411 3214 -339
<< psubdiffcont >>
rect -3201 -295 -3155 295
rect 3155 -295 3201 295
<< polysilicon >>
rect -2988 304 -2788 317
rect -2988 258 -2975 304
rect -2801 258 -2788 304
rect -2988 225 -2788 258
rect -2684 304 -2484 317
rect -2684 258 -2671 304
rect -2497 258 -2484 304
rect -2684 225 -2484 258
rect -2380 304 -2180 317
rect -2380 258 -2367 304
rect -2193 258 -2180 304
rect -2380 225 -2180 258
rect -2076 304 -1876 317
rect -2076 258 -2063 304
rect -1889 258 -1876 304
rect -2076 225 -1876 258
rect -1772 304 -1572 317
rect -1772 258 -1759 304
rect -1585 258 -1572 304
rect -1772 225 -1572 258
rect -1468 304 -1268 317
rect -1468 258 -1455 304
rect -1281 258 -1268 304
rect -1468 225 -1268 258
rect -1164 304 -964 317
rect -1164 258 -1151 304
rect -977 258 -964 304
rect -1164 225 -964 258
rect -860 304 -660 317
rect -860 258 -847 304
rect -673 258 -660 304
rect -860 225 -660 258
rect -556 304 -356 317
rect -556 258 -543 304
rect -369 258 -356 304
rect -556 225 -356 258
rect -252 304 -52 317
rect -252 258 -239 304
rect -65 258 -52 304
rect -252 225 -52 258
rect 52 304 252 317
rect 52 258 65 304
rect 239 258 252 304
rect 52 225 252 258
rect 356 304 556 317
rect 356 258 369 304
rect 543 258 556 304
rect 356 225 556 258
rect 660 304 860 317
rect 660 258 673 304
rect 847 258 860 304
rect 660 225 860 258
rect 964 304 1164 317
rect 964 258 977 304
rect 1151 258 1164 304
rect 964 225 1164 258
rect 1268 304 1468 317
rect 1268 258 1281 304
rect 1455 258 1468 304
rect 1268 225 1468 258
rect 1572 304 1772 317
rect 1572 258 1585 304
rect 1759 258 1772 304
rect 1572 225 1772 258
rect 1876 304 2076 317
rect 1876 258 1889 304
rect 2063 258 2076 304
rect 1876 225 2076 258
rect 2180 304 2380 317
rect 2180 258 2193 304
rect 2367 258 2380 304
rect 2180 225 2380 258
rect 2484 304 2684 317
rect 2484 258 2497 304
rect 2671 258 2684 304
rect 2484 225 2684 258
rect 2788 304 2988 317
rect 2788 258 2801 304
rect 2975 258 2988 304
rect 2788 225 2988 258
rect -2988 -258 -2788 -225
rect -2988 -304 -2975 -258
rect -2801 -304 -2788 -258
rect -2988 -317 -2788 -304
rect -2684 -258 -2484 -225
rect -2684 -304 -2671 -258
rect -2497 -304 -2484 -258
rect -2684 -317 -2484 -304
rect -2380 -258 -2180 -225
rect -2380 -304 -2367 -258
rect -2193 -304 -2180 -258
rect -2380 -317 -2180 -304
rect -2076 -258 -1876 -225
rect -2076 -304 -2063 -258
rect -1889 -304 -1876 -258
rect -2076 -317 -1876 -304
rect -1772 -258 -1572 -225
rect -1772 -304 -1759 -258
rect -1585 -304 -1572 -258
rect -1772 -317 -1572 -304
rect -1468 -258 -1268 -225
rect -1468 -304 -1455 -258
rect -1281 -304 -1268 -258
rect -1468 -317 -1268 -304
rect -1164 -258 -964 -225
rect -1164 -304 -1151 -258
rect -977 -304 -964 -258
rect -1164 -317 -964 -304
rect -860 -258 -660 -225
rect -860 -304 -847 -258
rect -673 -304 -660 -258
rect -860 -317 -660 -304
rect -556 -258 -356 -225
rect -556 -304 -543 -258
rect -369 -304 -356 -258
rect -556 -317 -356 -304
rect -252 -258 -52 -225
rect -252 -304 -239 -258
rect -65 -304 -52 -258
rect -252 -317 -52 -304
rect 52 -258 252 -225
rect 52 -304 65 -258
rect 239 -304 252 -258
rect 52 -317 252 -304
rect 356 -258 556 -225
rect 356 -304 369 -258
rect 543 -304 556 -258
rect 356 -317 556 -304
rect 660 -258 860 -225
rect 660 -304 673 -258
rect 847 -304 860 -258
rect 660 -317 860 -304
rect 964 -258 1164 -225
rect 964 -304 977 -258
rect 1151 -304 1164 -258
rect 964 -317 1164 -304
rect 1268 -258 1468 -225
rect 1268 -304 1281 -258
rect 1455 -304 1468 -258
rect 1268 -317 1468 -304
rect 1572 -258 1772 -225
rect 1572 -304 1585 -258
rect 1759 -304 1772 -258
rect 1572 -317 1772 -304
rect 1876 -258 2076 -225
rect 1876 -304 1889 -258
rect 2063 -304 2076 -258
rect 1876 -317 2076 -304
rect 2180 -258 2380 -225
rect 2180 -304 2193 -258
rect 2367 -304 2380 -258
rect 2180 -317 2380 -304
rect 2484 -258 2684 -225
rect 2484 -304 2497 -258
rect 2671 -304 2684 -258
rect 2484 -317 2684 -304
rect 2788 -258 2988 -225
rect 2788 -304 2801 -258
rect 2975 -304 2988 -258
rect 2788 -317 2988 -304
<< polycontact >>
rect -2975 258 -2801 304
rect -2671 258 -2497 304
rect -2367 258 -2193 304
rect -2063 258 -1889 304
rect -1759 258 -1585 304
rect -1455 258 -1281 304
rect -1151 258 -977 304
rect -847 258 -673 304
rect -543 258 -369 304
rect -239 258 -65 304
rect 65 258 239 304
rect 369 258 543 304
rect 673 258 847 304
rect 977 258 1151 304
rect 1281 258 1455 304
rect 1585 258 1759 304
rect 1889 258 2063 304
rect 2193 258 2367 304
rect 2497 258 2671 304
rect 2801 258 2975 304
rect -2975 -304 -2801 -258
rect -2671 -304 -2497 -258
rect -2367 -304 -2193 -258
rect -2063 -304 -1889 -258
rect -1759 -304 -1585 -258
rect -1455 -304 -1281 -258
rect -1151 -304 -977 -258
rect -847 -304 -673 -258
rect -543 -304 -369 -258
rect -239 -304 -65 -258
rect 65 -304 239 -258
rect 369 -304 543 -258
rect 673 -304 847 -258
rect 977 -304 1151 -258
rect 1281 -304 1455 -258
rect 1585 -304 1759 -258
rect 1889 -304 2063 -258
rect 2193 -304 2367 -258
rect 2497 -304 2671 -258
rect 2801 -304 2975 -258
<< metal1 >>
rect -3201 352 3201 398
rect -3201 295 -3155 352
rect -2986 258 -2975 304
rect -2801 258 -2790 304
rect -2682 258 -2671 304
rect -2497 258 -2486 304
rect -2378 258 -2367 304
rect -2193 258 -2182 304
rect -2074 258 -2063 304
rect -1889 258 -1878 304
rect -1770 258 -1759 304
rect -1585 258 -1574 304
rect -1466 258 -1455 304
rect -1281 258 -1270 304
rect -1162 258 -1151 304
rect -977 258 -966 304
rect -858 258 -847 304
rect -673 258 -662 304
rect -554 258 -543 304
rect -369 258 -358 304
rect -250 258 -239 304
rect -65 258 -54 304
rect 54 258 65 304
rect 239 258 250 304
rect 358 258 369 304
rect 543 258 554 304
rect 662 258 673 304
rect 847 258 858 304
rect 966 258 977 304
rect 1151 258 1162 304
rect 1270 258 1281 304
rect 1455 258 1466 304
rect 1574 258 1585 304
rect 1759 258 1770 304
rect 1878 258 1889 304
rect 2063 258 2074 304
rect 2182 258 2193 304
rect 2367 258 2378 304
rect 2486 258 2497 304
rect 2671 258 2682 304
rect 2790 258 2801 304
rect 2975 258 2986 304
rect 3155 295 3201 352
rect -3063 212 -3017 223
rect -3063 -223 -3017 -212
rect -2759 212 -2713 223
rect -2759 -223 -2713 -212
rect -2455 212 -2409 223
rect -2455 -223 -2409 -212
rect -2151 212 -2105 223
rect -2151 -223 -2105 -212
rect -1847 212 -1801 223
rect -1847 -223 -1801 -212
rect -1543 212 -1497 223
rect -1543 -223 -1497 -212
rect -1239 212 -1193 223
rect -1239 -223 -1193 -212
rect -935 212 -889 223
rect -935 -223 -889 -212
rect -631 212 -585 223
rect -631 -223 -585 -212
rect -327 212 -281 223
rect -327 -223 -281 -212
rect -23 212 23 223
rect -23 -223 23 -212
rect 281 212 327 223
rect 281 -223 327 -212
rect 585 212 631 223
rect 585 -223 631 -212
rect 889 212 935 223
rect 889 -223 935 -212
rect 1193 212 1239 223
rect 1193 -223 1239 -212
rect 1497 212 1543 223
rect 1497 -223 1543 -212
rect 1801 212 1847 223
rect 1801 -223 1847 -212
rect 2105 212 2151 223
rect 2105 -223 2151 -212
rect 2409 212 2455 223
rect 2409 -223 2455 -212
rect 2713 212 2759 223
rect 2713 -223 2759 -212
rect 3017 212 3063 223
rect 3017 -223 3063 -212
rect -3201 -352 -3155 -295
rect -2986 -304 -2975 -258
rect -2801 -304 -2790 -258
rect -2682 -304 -2671 -258
rect -2497 -304 -2486 -258
rect -2378 -304 -2367 -258
rect -2193 -304 -2182 -258
rect -2074 -304 -2063 -258
rect -1889 -304 -1878 -258
rect -1770 -304 -1759 -258
rect -1585 -304 -1574 -258
rect -1466 -304 -1455 -258
rect -1281 -304 -1270 -258
rect -1162 -304 -1151 -258
rect -977 -304 -966 -258
rect -858 -304 -847 -258
rect -673 -304 -662 -258
rect -554 -304 -543 -258
rect -369 -304 -358 -258
rect -250 -304 -239 -258
rect -65 -304 -54 -258
rect 54 -304 65 -258
rect 239 -304 250 -258
rect 358 -304 369 -258
rect 543 -304 554 -258
rect 662 -304 673 -258
rect 847 -304 858 -258
rect 966 -304 977 -258
rect 1151 -304 1162 -258
rect 1270 -304 1281 -258
rect 1455 -304 1466 -258
rect 1574 -304 1585 -258
rect 1759 -304 1770 -258
rect 1878 -304 1889 -258
rect 2063 -304 2074 -258
rect 2182 -304 2193 -258
rect 2367 -304 2378 -258
rect 2486 -304 2497 -258
rect 2671 -304 2682 -258
rect 2790 -304 2801 -258
rect 2975 -304 2986 -258
rect 3155 -352 3201 -295
rect -3201 -398 3201 -352
<< properties >>
string FIXED_BBOX -3178 -375 3178 375
string gencell nfet_03v3
string library gf180mcu
string parameters w 2.25 l 1.0 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
