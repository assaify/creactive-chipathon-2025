magic
tech gf180mcuD
magscale 1 10
timestamp 1755278675
<< mimcap >>
rect -12883 5640 -10883 5720
rect -12883 3800 -12803 5640
rect -10963 3800 -10883 5640
rect -12883 3720 -10883 3800
rect -10269 5640 -8269 5720
rect -10269 3800 -10189 5640
rect -8349 3800 -8269 5640
rect -10269 3720 -8269 3800
rect -7655 5640 -5655 5720
rect -7655 3800 -7575 5640
rect -5735 3800 -5655 5640
rect -7655 3720 -5655 3800
rect -5041 5640 -3041 5720
rect -5041 3800 -4961 5640
rect -3121 3800 -3041 5640
rect -5041 3720 -3041 3800
rect -2427 5640 -427 5720
rect -2427 3800 -2347 5640
rect -507 3800 -427 5640
rect -2427 3720 -427 3800
rect 187 5640 2187 5720
rect 187 3800 267 5640
rect 2107 3800 2187 5640
rect 187 3720 2187 3800
rect 2801 5640 4801 5720
rect 2801 3800 2881 5640
rect 4721 3800 4801 5640
rect 2801 3720 4801 3800
rect 5415 5640 7415 5720
rect 5415 3800 5495 5640
rect 7335 3800 7415 5640
rect 5415 3720 7415 3800
rect 8029 5640 10029 5720
rect 8029 3800 8109 5640
rect 9949 3800 10029 5640
rect 8029 3720 10029 3800
rect 10643 5640 12643 5720
rect 10643 3800 10723 5640
rect 12563 3800 12643 5640
rect 10643 3720 12643 3800
rect -12883 3280 -10883 3360
rect -12883 1440 -12803 3280
rect -10963 1440 -10883 3280
rect -12883 1360 -10883 1440
rect -10269 3280 -8269 3360
rect -10269 1440 -10189 3280
rect -8349 1440 -8269 3280
rect -10269 1360 -8269 1440
rect -7655 3280 -5655 3360
rect -7655 1440 -7575 3280
rect -5735 1440 -5655 3280
rect -7655 1360 -5655 1440
rect -5041 3280 -3041 3360
rect -5041 1440 -4961 3280
rect -3121 1440 -3041 3280
rect -5041 1360 -3041 1440
rect -2427 3280 -427 3360
rect -2427 1440 -2347 3280
rect -507 1440 -427 3280
rect -2427 1360 -427 1440
rect 187 3280 2187 3360
rect 187 1440 267 3280
rect 2107 1440 2187 3280
rect 187 1360 2187 1440
rect 2801 3280 4801 3360
rect 2801 1440 2881 3280
rect 4721 1440 4801 3280
rect 2801 1360 4801 1440
rect 5415 3280 7415 3360
rect 5415 1440 5495 3280
rect 7335 1440 7415 3280
rect 5415 1360 7415 1440
rect 8029 3280 10029 3360
rect 8029 1440 8109 3280
rect 9949 1440 10029 3280
rect 8029 1360 10029 1440
rect 10643 3280 12643 3360
rect 10643 1440 10723 3280
rect 12563 1440 12643 3280
rect 10643 1360 12643 1440
rect -12883 920 -10883 1000
rect -12883 -920 -12803 920
rect -10963 -920 -10883 920
rect -12883 -1000 -10883 -920
rect -10269 920 -8269 1000
rect -10269 -920 -10189 920
rect -8349 -920 -8269 920
rect -10269 -1000 -8269 -920
rect -7655 920 -5655 1000
rect -7655 -920 -7575 920
rect -5735 -920 -5655 920
rect -7655 -1000 -5655 -920
rect -5041 920 -3041 1000
rect -5041 -920 -4961 920
rect -3121 -920 -3041 920
rect -5041 -1000 -3041 -920
rect -2427 920 -427 1000
rect -2427 -920 -2347 920
rect -507 -920 -427 920
rect -2427 -1000 -427 -920
rect 187 920 2187 1000
rect 187 -920 267 920
rect 2107 -920 2187 920
rect 187 -1000 2187 -920
rect 2801 920 4801 1000
rect 2801 -920 2881 920
rect 4721 -920 4801 920
rect 2801 -1000 4801 -920
rect 5415 920 7415 1000
rect 5415 -920 5495 920
rect 7335 -920 7415 920
rect 5415 -1000 7415 -920
rect 8029 920 10029 1000
rect 8029 -920 8109 920
rect 9949 -920 10029 920
rect 8029 -1000 10029 -920
rect 10643 920 12643 1000
rect 10643 -920 10723 920
rect 12563 -920 12643 920
rect 10643 -1000 12643 -920
rect -12883 -1440 -10883 -1360
rect -12883 -3280 -12803 -1440
rect -10963 -3280 -10883 -1440
rect -12883 -3360 -10883 -3280
rect -10269 -1440 -8269 -1360
rect -10269 -3280 -10189 -1440
rect -8349 -3280 -8269 -1440
rect -10269 -3360 -8269 -3280
rect -7655 -1440 -5655 -1360
rect -7655 -3280 -7575 -1440
rect -5735 -3280 -5655 -1440
rect -7655 -3360 -5655 -3280
rect -5041 -1440 -3041 -1360
rect -5041 -3280 -4961 -1440
rect -3121 -3280 -3041 -1440
rect -5041 -3360 -3041 -3280
rect -2427 -1440 -427 -1360
rect -2427 -3280 -2347 -1440
rect -507 -3280 -427 -1440
rect -2427 -3360 -427 -3280
rect 187 -1440 2187 -1360
rect 187 -3280 267 -1440
rect 2107 -3280 2187 -1440
rect 187 -3360 2187 -3280
rect 2801 -1440 4801 -1360
rect 2801 -3280 2881 -1440
rect 4721 -3280 4801 -1440
rect 2801 -3360 4801 -3280
rect 5415 -1440 7415 -1360
rect 5415 -3280 5495 -1440
rect 7335 -3280 7415 -1440
rect 5415 -3360 7415 -3280
rect 8029 -1440 10029 -1360
rect 8029 -3280 8109 -1440
rect 9949 -3280 10029 -1440
rect 8029 -3360 10029 -3280
rect 10643 -1440 12643 -1360
rect 10643 -3280 10723 -1440
rect 12563 -3280 12643 -1440
rect 10643 -3360 12643 -3280
rect -12883 -3800 -10883 -3720
rect -12883 -5640 -12803 -3800
rect -10963 -5640 -10883 -3800
rect -12883 -5720 -10883 -5640
rect -10269 -3800 -8269 -3720
rect -10269 -5640 -10189 -3800
rect -8349 -5640 -8269 -3800
rect -10269 -5720 -8269 -5640
rect -7655 -3800 -5655 -3720
rect -7655 -5640 -7575 -3800
rect -5735 -5640 -5655 -3800
rect -7655 -5720 -5655 -5640
rect -5041 -3800 -3041 -3720
rect -5041 -5640 -4961 -3800
rect -3121 -5640 -3041 -3800
rect -5041 -5720 -3041 -5640
rect -2427 -3800 -427 -3720
rect -2427 -5640 -2347 -3800
rect -507 -5640 -427 -3800
rect -2427 -5720 -427 -5640
rect 187 -3800 2187 -3720
rect 187 -5640 267 -3800
rect 2107 -5640 2187 -3800
rect 187 -5720 2187 -5640
rect 2801 -3800 4801 -3720
rect 2801 -5640 2881 -3800
rect 4721 -5640 4801 -3800
rect 2801 -5720 4801 -5640
rect 5415 -3800 7415 -3720
rect 5415 -5640 5495 -3800
rect 7335 -5640 7415 -3800
rect 5415 -5720 7415 -5640
rect 8029 -3800 10029 -3720
rect 8029 -5640 8109 -3800
rect 9949 -5640 10029 -3800
rect 8029 -5720 10029 -5640
rect 10643 -3800 12643 -3720
rect 10643 -5640 10723 -3800
rect 12563 -5640 12643 -3800
rect 10643 -5720 12643 -5640
<< mimcapcontact >>
rect -12803 3800 -10963 5640
rect -10189 3800 -8349 5640
rect -7575 3800 -5735 5640
rect -4961 3800 -3121 5640
rect -2347 3800 -507 5640
rect 267 3800 2107 5640
rect 2881 3800 4721 5640
rect 5495 3800 7335 5640
rect 8109 3800 9949 5640
rect 10723 3800 12563 5640
rect -12803 1440 -10963 3280
rect -10189 1440 -8349 3280
rect -7575 1440 -5735 3280
rect -4961 1440 -3121 3280
rect -2347 1440 -507 3280
rect 267 1440 2107 3280
rect 2881 1440 4721 3280
rect 5495 1440 7335 3280
rect 8109 1440 9949 3280
rect 10723 1440 12563 3280
rect -12803 -920 -10963 920
rect -10189 -920 -8349 920
rect -7575 -920 -5735 920
rect -4961 -920 -3121 920
rect -2347 -920 -507 920
rect 267 -920 2107 920
rect 2881 -920 4721 920
rect 5495 -920 7335 920
rect 8109 -920 9949 920
rect 10723 -920 12563 920
rect -12803 -3280 -10963 -1440
rect -10189 -3280 -8349 -1440
rect -7575 -3280 -5735 -1440
rect -4961 -3280 -3121 -1440
rect -2347 -3280 -507 -1440
rect 267 -3280 2107 -1440
rect 2881 -3280 4721 -1440
rect 5495 -3280 7335 -1440
rect 8109 -3280 9949 -1440
rect 10723 -3280 12563 -1440
rect -12803 -5640 -10963 -3800
rect -10189 -5640 -8349 -3800
rect -7575 -5640 -5735 -3800
rect -4961 -5640 -3121 -3800
rect -2347 -5640 -507 -3800
rect 267 -5640 2107 -3800
rect 2881 -5640 4721 -3800
rect 5495 -5640 7335 -3800
rect 8109 -5640 9949 -3800
rect 10723 -5640 12563 -3800
<< metal4 >>
rect -13003 5773 -10523 5840
rect -13003 5720 -10673 5773
rect -13003 3720 -12883 5720
rect -10883 3720 -10673 5720
rect -13003 3667 -10673 3720
rect -10585 3667 -10523 5773
rect -13003 3600 -10523 3667
rect -10389 5773 -7909 5840
rect -10389 5720 -8059 5773
rect -10389 3720 -10269 5720
rect -8269 3720 -8059 5720
rect -10389 3667 -8059 3720
rect -7971 3667 -7909 5773
rect -10389 3600 -7909 3667
rect -7775 5773 -5295 5840
rect -7775 5720 -5445 5773
rect -7775 3720 -7655 5720
rect -5655 3720 -5445 5720
rect -7775 3667 -5445 3720
rect -5357 3667 -5295 5773
rect -7775 3600 -5295 3667
rect -5161 5773 -2681 5840
rect -5161 5720 -2831 5773
rect -5161 3720 -5041 5720
rect -3041 3720 -2831 5720
rect -5161 3667 -2831 3720
rect -2743 3667 -2681 5773
rect -5161 3600 -2681 3667
rect -2547 5773 -67 5840
rect -2547 5720 -217 5773
rect -2547 3720 -2427 5720
rect -427 3720 -217 5720
rect -2547 3667 -217 3720
rect -129 3667 -67 5773
rect -2547 3600 -67 3667
rect 67 5773 2547 5840
rect 67 5720 2397 5773
rect 67 3720 187 5720
rect 2187 3720 2397 5720
rect 67 3667 2397 3720
rect 2485 3667 2547 5773
rect 67 3600 2547 3667
rect 2681 5773 5161 5840
rect 2681 5720 5011 5773
rect 2681 3720 2801 5720
rect 4801 3720 5011 5720
rect 2681 3667 5011 3720
rect 5099 3667 5161 5773
rect 2681 3600 5161 3667
rect 5295 5773 7775 5840
rect 5295 5720 7625 5773
rect 5295 3720 5415 5720
rect 7415 3720 7625 5720
rect 5295 3667 7625 3720
rect 7713 3667 7775 5773
rect 5295 3600 7775 3667
rect 7909 5773 10389 5840
rect 7909 5720 10239 5773
rect 7909 3720 8029 5720
rect 10029 3720 10239 5720
rect 7909 3667 10239 3720
rect 10327 3667 10389 5773
rect 7909 3600 10389 3667
rect 10523 5773 13003 5840
rect 10523 5720 12853 5773
rect 10523 3720 10643 5720
rect 12643 3720 12853 5720
rect 10523 3667 12853 3720
rect 12941 3667 13003 5773
rect 10523 3600 13003 3667
rect -13003 3413 -10523 3480
rect -13003 3360 -10673 3413
rect -13003 1360 -12883 3360
rect -10883 1360 -10673 3360
rect -13003 1307 -10673 1360
rect -10585 1307 -10523 3413
rect -13003 1240 -10523 1307
rect -10389 3413 -7909 3480
rect -10389 3360 -8059 3413
rect -10389 1360 -10269 3360
rect -8269 1360 -8059 3360
rect -10389 1307 -8059 1360
rect -7971 1307 -7909 3413
rect -10389 1240 -7909 1307
rect -7775 3413 -5295 3480
rect -7775 3360 -5445 3413
rect -7775 1360 -7655 3360
rect -5655 1360 -5445 3360
rect -7775 1307 -5445 1360
rect -5357 1307 -5295 3413
rect -7775 1240 -5295 1307
rect -5161 3413 -2681 3480
rect -5161 3360 -2831 3413
rect -5161 1360 -5041 3360
rect -3041 1360 -2831 3360
rect -5161 1307 -2831 1360
rect -2743 1307 -2681 3413
rect -5161 1240 -2681 1307
rect -2547 3413 -67 3480
rect -2547 3360 -217 3413
rect -2547 1360 -2427 3360
rect -427 1360 -217 3360
rect -2547 1307 -217 1360
rect -129 1307 -67 3413
rect -2547 1240 -67 1307
rect 67 3413 2547 3480
rect 67 3360 2397 3413
rect 67 1360 187 3360
rect 2187 1360 2397 3360
rect 67 1307 2397 1360
rect 2485 1307 2547 3413
rect 67 1240 2547 1307
rect 2681 3413 5161 3480
rect 2681 3360 5011 3413
rect 2681 1360 2801 3360
rect 4801 1360 5011 3360
rect 2681 1307 5011 1360
rect 5099 1307 5161 3413
rect 2681 1240 5161 1307
rect 5295 3413 7775 3480
rect 5295 3360 7625 3413
rect 5295 1360 5415 3360
rect 7415 1360 7625 3360
rect 5295 1307 7625 1360
rect 7713 1307 7775 3413
rect 5295 1240 7775 1307
rect 7909 3413 10389 3480
rect 7909 3360 10239 3413
rect 7909 1360 8029 3360
rect 10029 1360 10239 3360
rect 7909 1307 10239 1360
rect 10327 1307 10389 3413
rect 7909 1240 10389 1307
rect 10523 3413 13003 3480
rect 10523 3360 12853 3413
rect 10523 1360 10643 3360
rect 12643 1360 12853 3360
rect 10523 1307 12853 1360
rect 12941 1307 13003 3413
rect 10523 1240 13003 1307
rect -13003 1053 -10523 1120
rect -13003 1000 -10673 1053
rect -13003 -1000 -12883 1000
rect -10883 -1000 -10673 1000
rect -13003 -1053 -10673 -1000
rect -10585 -1053 -10523 1053
rect -13003 -1120 -10523 -1053
rect -10389 1053 -7909 1120
rect -10389 1000 -8059 1053
rect -10389 -1000 -10269 1000
rect -8269 -1000 -8059 1000
rect -10389 -1053 -8059 -1000
rect -7971 -1053 -7909 1053
rect -10389 -1120 -7909 -1053
rect -7775 1053 -5295 1120
rect -7775 1000 -5445 1053
rect -7775 -1000 -7655 1000
rect -5655 -1000 -5445 1000
rect -7775 -1053 -5445 -1000
rect -5357 -1053 -5295 1053
rect -7775 -1120 -5295 -1053
rect -5161 1053 -2681 1120
rect -5161 1000 -2831 1053
rect -5161 -1000 -5041 1000
rect -3041 -1000 -2831 1000
rect -5161 -1053 -2831 -1000
rect -2743 -1053 -2681 1053
rect -5161 -1120 -2681 -1053
rect -2547 1053 -67 1120
rect -2547 1000 -217 1053
rect -2547 -1000 -2427 1000
rect -427 -1000 -217 1000
rect -2547 -1053 -217 -1000
rect -129 -1053 -67 1053
rect -2547 -1120 -67 -1053
rect 67 1053 2547 1120
rect 67 1000 2397 1053
rect 67 -1000 187 1000
rect 2187 -1000 2397 1000
rect 67 -1053 2397 -1000
rect 2485 -1053 2547 1053
rect 67 -1120 2547 -1053
rect 2681 1053 5161 1120
rect 2681 1000 5011 1053
rect 2681 -1000 2801 1000
rect 4801 -1000 5011 1000
rect 2681 -1053 5011 -1000
rect 5099 -1053 5161 1053
rect 2681 -1120 5161 -1053
rect 5295 1053 7775 1120
rect 5295 1000 7625 1053
rect 5295 -1000 5415 1000
rect 7415 -1000 7625 1000
rect 5295 -1053 7625 -1000
rect 7713 -1053 7775 1053
rect 5295 -1120 7775 -1053
rect 7909 1053 10389 1120
rect 7909 1000 10239 1053
rect 7909 -1000 8029 1000
rect 10029 -1000 10239 1000
rect 7909 -1053 10239 -1000
rect 10327 -1053 10389 1053
rect 7909 -1120 10389 -1053
rect 10523 1053 13003 1120
rect 10523 1000 12853 1053
rect 10523 -1000 10643 1000
rect 12643 -1000 12853 1000
rect 10523 -1053 12853 -1000
rect 12941 -1053 13003 1053
rect 10523 -1120 13003 -1053
rect -13003 -1307 -10523 -1240
rect -13003 -1360 -10673 -1307
rect -13003 -3360 -12883 -1360
rect -10883 -3360 -10673 -1360
rect -13003 -3413 -10673 -3360
rect -10585 -3413 -10523 -1307
rect -13003 -3480 -10523 -3413
rect -10389 -1307 -7909 -1240
rect -10389 -1360 -8059 -1307
rect -10389 -3360 -10269 -1360
rect -8269 -3360 -8059 -1360
rect -10389 -3413 -8059 -3360
rect -7971 -3413 -7909 -1307
rect -10389 -3480 -7909 -3413
rect -7775 -1307 -5295 -1240
rect -7775 -1360 -5445 -1307
rect -7775 -3360 -7655 -1360
rect -5655 -3360 -5445 -1360
rect -7775 -3413 -5445 -3360
rect -5357 -3413 -5295 -1307
rect -7775 -3480 -5295 -3413
rect -5161 -1307 -2681 -1240
rect -5161 -1360 -2831 -1307
rect -5161 -3360 -5041 -1360
rect -3041 -3360 -2831 -1360
rect -5161 -3413 -2831 -3360
rect -2743 -3413 -2681 -1307
rect -5161 -3480 -2681 -3413
rect -2547 -1307 -67 -1240
rect -2547 -1360 -217 -1307
rect -2547 -3360 -2427 -1360
rect -427 -3360 -217 -1360
rect -2547 -3413 -217 -3360
rect -129 -3413 -67 -1307
rect -2547 -3480 -67 -3413
rect 67 -1307 2547 -1240
rect 67 -1360 2397 -1307
rect 67 -3360 187 -1360
rect 2187 -3360 2397 -1360
rect 67 -3413 2397 -3360
rect 2485 -3413 2547 -1307
rect 67 -3480 2547 -3413
rect 2681 -1307 5161 -1240
rect 2681 -1360 5011 -1307
rect 2681 -3360 2801 -1360
rect 4801 -3360 5011 -1360
rect 2681 -3413 5011 -3360
rect 5099 -3413 5161 -1307
rect 2681 -3480 5161 -3413
rect 5295 -1307 7775 -1240
rect 5295 -1360 7625 -1307
rect 5295 -3360 5415 -1360
rect 7415 -3360 7625 -1360
rect 5295 -3413 7625 -3360
rect 7713 -3413 7775 -1307
rect 5295 -3480 7775 -3413
rect 7909 -1307 10389 -1240
rect 7909 -1360 10239 -1307
rect 7909 -3360 8029 -1360
rect 10029 -3360 10239 -1360
rect 7909 -3413 10239 -3360
rect 10327 -3413 10389 -1307
rect 7909 -3480 10389 -3413
rect 10523 -1307 13003 -1240
rect 10523 -1360 12853 -1307
rect 10523 -3360 10643 -1360
rect 12643 -3360 12853 -1360
rect 10523 -3413 12853 -3360
rect 12941 -3413 13003 -1307
rect 10523 -3480 13003 -3413
rect -13003 -3667 -10523 -3600
rect -13003 -3720 -10673 -3667
rect -13003 -5720 -12883 -3720
rect -10883 -5720 -10673 -3720
rect -13003 -5773 -10673 -5720
rect -10585 -5773 -10523 -3667
rect -13003 -5840 -10523 -5773
rect -10389 -3667 -7909 -3600
rect -10389 -3720 -8059 -3667
rect -10389 -5720 -10269 -3720
rect -8269 -5720 -8059 -3720
rect -10389 -5773 -8059 -5720
rect -7971 -5773 -7909 -3667
rect -10389 -5840 -7909 -5773
rect -7775 -3667 -5295 -3600
rect -7775 -3720 -5445 -3667
rect -7775 -5720 -7655 -3720
rect -5655 -5720 -5445 -3720
rect -7775 -5773 -5445 -5720
rect -5357 -5773 -5295 -3667
rect -7775 -5840 -5295 -5773
rect -5161 -3667 -2681 -3600
rect -5161 -3720 -2831 -3667
rect -5161 -5720 -5041 -3720
rect -3041 -5720 -2831 -3720
rect -5161 -5773 -2831 -5720
rect -2743 -5773 -2681 -3667
rect -5161 -5840 -2681 -5773
rect -2547 -3667 -67 -3600
rect -2547 -3720 -217 -3667
rect -2547 -5720 -2427 -3720
rect -427 -5720 -217 -3720
rect -2547 -5773 -217 -5720
rect -129 -5773 -67 -3667
rect -2547 -5840 -67 -5773
rect 67 -3667 2547 -3600
rect 67 -3720 2397 -3667
rect 67 -5720 187 -3720
rect 2187 -5720 2397 -3720
rect 67 -5773 2397 -5720
rect 2485 -5773 2547 -3667
rect 67 -5840 2547 -5773
rect 2681 -3667 5161 -3600
rect 2681 -3720 5011 -3667
rect 2681 -5720 2801 -3720
rect 4801 -5720 5011 -3720
rect 2681 -5773 5011 -5720
rect 5099 -5773 5161 -3667
rect 2681 -5840 5161 -5773
rect 5295 -3667 7775 -3600
rect 5295 -3720 7625 -3667
rect 5295 -5720 5415 -3720
rect 7415 -5720 7625 -3720
rect 5295 -5773 7625 -5720
rect 7713 -5773 7775 -3667
rect 5295 -5840 7775 -5773
rect 7909 -3667 10389 -3600
rect 7909 -3720 10239 -3667
rect 7909 -5720 8029 -3720
rect 10029 -5720 10239 -3720
rect 7909 -5773 10239 -5720
rect 10327 -5773 10389 -3667
rect 7909 -5840 10389 -5773
rect 10523 -3667 13003 -3600
rect 10523 -3720 12853 -3667
rect 10523 -5720 10643 -3720
rect 12643 -5720 12853 -3720
rect 10523 -5773 12853 -5720
rect 12941 -5773 13003 -3667
rect 10523 -5840 13003 -5773
<< via4 >>
rect -10673 3667 -10585 5773
rect -8059 3667 -7971 5773
rect -5445 3667 -5357 5773
rect -2831 3667 -2743 5773
rect -217 3667 -129 5773
rect 2397 3667 2485 5773
rect 5011 3667 5099 5773
rect 7625 3667 7713 5773
rect 10239 3667 10327 5773
rect 12853 3667 12941 5773
rect -10673 1307 -10585 3413
rect -8059 1307 -7971 3413
rect -5445 1307 -5357 3413
rect -2831 1307 -2743 3413
rect -217 1307 -129 3413
rect 2397 1307 2485 3413
rect 5011 1307 5099 3413
rect 7625 1307 7713 3413
rect 10239 1307 10327 3413
rect 12853 1307 12941 3413
rect -10673 -1053 -10585 1053
rect -8059 -1053 -7971 1053
rect -5445 -1053 -5357 1053
rect -2831 -1053 -2743 1053
rect -217 -1053 -129 1053
rect 2397 -1053 2485 1053
rect 5011 -1053 5099 1053
rect 7625 -1053 7713 1053
rect 10239 -1053 10327 1053
rect 12853 -1053 12941 1053
rect -10673 -3413 -10585 -1307
rect -8059 -3413 -7971 -1307
rect -5445 -3413 -5357 -1307
rect -2831 -3413 -2743 -1307
rect -217 -3413 -129 -1307
rect 2397 -3413 2485 -1307
rect 5011 -3413 5099 -1307
rect 7625 -3413 7713 -1307
rect 10239 -3413 10327 -1307
rect 12853 -3413 12941 -1307
rect -10673 -5773 -10585 -3667
rect -8059 -5773 -7971 -3667
rect -5445 -5773 -5357 -3667
rect -2831 -5773 -2743 -3667
rect -217 -5773 -129 -3667
rect 2397 -5773 2485 -3667
rect 5011 -5773 5099 -3667
rect 7625 -5773 7713 -3667
rect 10239 -5773 10327 -3667
rect 12853 -5773 12941 -3667
<< metal5 >>
rect -11989 5640 -11777 5900
rect -10735 5773 -10523 5900
rect -11989 3280 -11777 3800
rect -10735 3667 -10673 5773
rect -10585 3667 -10523 5773
rect -9375 5640 -9163 5900
rect -8121 5773 -7909 5900
rect -10735 3413 -10523 3667
rect -11989 920 -11777 1440
rect -10735 1307 -10673 3413
rect -10585 1307 -10523 3413
rect -9375 3280 -9163 3800
rect -8121 3667 -8059 5773
rect -7971 3667 -7909 5773
rect -6761 5640 -6549 5900
rect -5507 5773 -5295 5900
rect -8121 3413 -7909 3667
rect -10735 1053 -10523 1307
rect -11989 -1440 -11777 -920
rect -10735 -1053 -10673 1053
rect -10585 -1053 -10523 1053
rect -9375 920 -9163 1440
rect -8121 1307 -8059 3413
rect -7971 1307 -7909 3413
rect -6761 3280 -6549 3800
rect -5507 3667 -5445 5773
rect -5357 3667 -5295 5773
rect -4147 5640 -3935 5900
rect -2893 5773 -2681 5900
rect -5507 3413 -5295 3667
rect -8121 1053 -7909 1307
rect -10735 -1307 -10523 -1053
rect -11989 -3800 -11777 -3280
rect -10735 -3413 -10673 -1307
rect -10585 -3413 -10523 -1307
rect -9375 -1440 -9163 -920
rect -8121 -1053 -8059 1053
rect -7971 -1053 -7909 1053
rect -6761 920 -6549 1440
rect -5507 1307 -5445 3413
rect -5357 1307 -5295 3413
rect -4147 3280 -3935 3800
rect -2893 3667 -2831 5773
rect -2743 3667 -2681 5773
rect -1533 5640 -1321 5900
rect -279 5773 -67 5900
rect -2893 3413 -2681 3667
rect -5507 1053 -5295 1307
rect -8121 -1307 -7909 -1053
rect -10735 -3667 -10523 -3413
rect -11989 -5900 -11777 -5640
rect -10735 -5773 -10673 -3667
rect -10585 -5773 -10523 -3667
rect -9375 -3800 -9163 -3280
rect -8121 -3413 -8059 -1307
rect -7971 -3413 -7909 -1307
rect -6761 -1440 -6549 -920
rect -5507 -1053 -5445 1053
rect -5357 -1053 -5295 1053
rect -4147 920 -3935 1440
rect -2893 1307 -2831 3413
rect -2743 1307 -2681 3413
rect -1533 3280 -1321 3800
rect -279 3667 -217 5773
rect -129 3667 -67 5773
rect 1081 5640 1293 5900
rect 2335 5773 2547 5900
rect -279 3413 -67 3667
rect -2893 1053 -2681 1307
rect -5507 -1307 -5295 -1053
rect -8121 -3667 -7909 -3413
rect -10735 -5900 -10523 -5773
rect -9375 -5900 -9163 -5640
rect -8121 -5773 -8059 -3667
rect -7971 -5773 -7909 -3667
rect -6761 -3800 -6549 -3280
rect -5507 -3413 -5445 -1307
rect -5357 -3413 -5295 -1307
rect -4147 -1440 -3935 -920
rect -2893 -1053 -2831 1053
rect -2743 -1053 -2681 1053
rect -1533 920 -1321 1440
rect -279 1307 -217 3413
rect -129 1307 -67 3413
rect 1081 3280 1293 3800
rect 2335 3667 2397 5773
rect 2485 3667 2547 5773
rect 3695 5640 3907 5900
rect 4949 5773 5161 5900
rect 2335 3413 2547 3667
rect -279 1053 -67 1307
rect -2893 -1307 -2681 -1053
rect -5507 -3667 -5295 -3413
rect -8121 -5900 -7909 -5773
rect -6761 -5900 -6549 -5640
rect -5507 -5773 -5445 -3667
rect -5357 -5773 -5295 -3667
rect -4147 -3800 -3935 -3280
rect -2893 -3413 -2831 -1307
rect -2743 -3413 -2681 -1307
rect -1533 -1440 -1321 -920
rect -279 -1053 -217 1053
rect -129 -1053 -67 1053
rect 1081 920 1293 1440
rect 2335 1307 2397 3413
rect 2485 1307 2547 3413
rect 3695 3280 3907 3800
rect 4949 3667 5011 5773
rect 5099 3667 5161 5773
rect 6309 5640 6521 5900
rect 7563 5773 7775 5900
rect 4949 3413 5161 3667
rect 2335 1053 2547 1307
rect -279 -1307 -67 -1053
rect -2893 -3667 -2681 -3413
rect -5507 -5900 -5295 -5773
rect -4147 -5900 -3935 -5640
rect -2893 -5773 -2831 -3667
rect -2743 -5773 -2681 -3667
rect -1533 -3800 -1321 -3280
rect -279 -3413 -217 -1307
rect -129 -3413 -67 -1307
rect 1081 -1440 1293 -920
rect 2335 -1053 2397 1053
rect 2485 -1053 2547 1053
rect 3695 920 3907 1440
rect 4949 1307 5011 3413
rect 5099 1307 5161 3413
rect 6309 3280 6521 3800
rect 7563 3667 7625 5773
rect 7713 3667 7775 5773
rect 8923 5640 9135 5900
rect 10177 5773 10389 5900
rect 7563 3413 7775 3667
rect 4949 1053 5161 1307
rect 2335 -1307 2547 -1053
rect -279 -3667 -67 -3413
rect -2893 -5900 -2681 -5773
rect -1533 -5900 -1321 -5640
rect -279 -5773 -217 -3667
rect -129 -5773 -67 -3667
rect 1081 -3800 1293 -3280
rect 2335 -3413 2397 -1307
rect 2485 -3413 2547 -1307
rect 3695 -1440 3907 -920
rect 4949 -1053 5011 1053
rect 5099 -1053 5161 1053
rect 6309 920 6521 1440
rect 7563 1307 7625 3413
rect 7713 1307 7775 3413
rect 8923 3280 9135 3800
rect 10177 3667 10239 5773
rect 10327 3667 10389 5773
rect 11537 5640 11749 5900
rect 12791 5773 13003 5900
rect 10177 3413 10389 3667
rect 7563 1053 7775 1307
rect 4949 -1307 5161 -1053
rect 2335 -3667 2547 -3413
rect -279 -5900 -67 -5773
rect 1081 -5900 1293 -5640
rect 2335 -5773 2397 -3667
rect 2485 -5773 2547 -3667
rect 3695 -3800 3907 -3280
rect 4949 -3413 5011 -1307
rect 5099 -3413 5161 -1307
rect 6309 -1440 6521 -920
rect 7563 -1053 7625 1053
rect 7713 -1053 7775 1053
rect 8923 920 9135 1440
rect 10177 1307 10239 3413
rect 10327 1307 10389 3413
rect 11537 3280 11749 3800
rect 12791 3667 12853 5773
rect 12941 3667 13003 5773
rect 12791 3413 13003 3667
rect 10177 1053 10389 1307
rect 7563 -1307 7775 -1053
rect 4949 -3667 5161 -3413
rect 2335 -5900 2547 -5773
rect 3695 -5900 3907 -5640
rect 4949 -5773 5011 -3667
rect 5099 -5773 5161 -3667
rect 6309 -3800 6521 -3280
rect 7563 -3413 7625 -1307
rect 7713 -3413 7775 -1307
rect 8923 -1440 9135 -920
rect 10177 -1053 10239 1053
rect 10327 -1053 10389 1053
rect 11537 920 11749 1440
rect 12791 1307 12853 3413
rect 12941 1307 13003 3413
rect 12791 1053 13003 1307
rect 10177 -1307 10389 -1053
rect 7563 -3667 7775 -3413
rect 4949 -5900 5161 -5773
rect 6309 -5900 6521 -5640
rect 7563 -5773 7625 -3667
rect 7713 -5773 7775 -3667
rect 8923 -3800 9135 -3280
rect 10177 -3413 10239 -1307
rect 10327 -3413 10389 -1307
rect 11537 -1440 11749 -920
rect 12791 -1053 12853 1053
rect 12941 -1053 13003 1053
rect 12791 -1307 13003 -1053
rect 10177 -3667 10389 -3413
rect 7563 -5900 7775 -5773
rect 8923 -5900 9135 -5640
rect 10177 -5773 10239 -3667
rect 10327 -5773 10389 -3667
rect 11537 -3800 11749 -3280
rect 12791 -3413 12853 -1307
rect 12941 -3413 13003 -1307
rect 12791 -3667 13003 -3413
rect 10177 -5900 10389 -5773
rect 11537 -5900 11749 -5640
rect 12791 -5773 12853 -3667
rect 12941 -5773 13003 -3667
rect 12791 -5900 13003 -5773
<< properties >>
string FIXED_BBOX 10523 3600 12763 5840
string gencell cap_mim_2p0fF
string library gf180mcu
string parameters w 10 l 10 val 3.3k carea 25.00 cperi 20.00 class capacitor nx 10 ny 5 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 1 tconnect 1
<< end >>
