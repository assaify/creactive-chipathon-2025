magic
tech gf180mcuD
magscale 1 10
timestamp 1758305657
<< psubdiff >>
rect -1321 1642 12391 1669
rect -1321 1596 -1169 1642
rect 12239 1596 12391 1642
rect -1321 1569 12391 1596
rect -1321 1444 -1221 1569
rect -1321 -1050 -1294 1444
rect -1248 -1050 -1221 1444
rect -1321 -1175 -1221 -1050
rect 12291 1444 12391 1569
rect 12291 -1050 12318 1444
rect 12364 -1050 12391 1444
rect 12291 -1175 12391 -1050
rect -1321 -1202 12391 -1175
rect -1321 -1248 -1169 -1202
rect 12239 -1248 12391 -1202
rect -1321 -1275 12391 -1248
<< psubdiffcont >>
rect -1169 1596 12239 1642
rect -1294 -1050 -1248 1444
rect 12318 -1050 12364 1444
rect -1169 -1248 12239 -1202
<< metal1 >>
rect -1357 1645 12427 1705
rect -1357 1642 -801 1645
rect -749 1642 2057 1645
rect 2109 1642 2453 1645
rect 2505 1642 5311 1645
rect 5363 1642 5707 1645
rect 5759 1642 8565 1645
rect 8617 1642 8961 1645
rect 9013 1642 11819 1645
rect 11871 1642 12427 1645
rect -1357 1596 -1169 1642
rect 12239 1596 12427 1642
rect -1357 1593 -801 1596
rect -749 1593 2057 1596
rect 2109 1593 2453 1596
rect 2505 1593 5311 1596
rect 5363 1593 5707 1596
rect 5759 1593 8565 1596
rect 8617 1593 8961 1596
rect 9013 1593 11819 1596
rect 11871 1593 12427 1596
rect -1357 1533 12427 1593
rect -1357 1444 -1185 1533
rect -1357 -1050 -1294 1444
rect -1248 -1050 -1185 1444
rect -965 1449 12142 1473
rect -965 1397 2321 1449
rect 2373 1397 8829 1449
rect 8881 1397 12142 1449
rect -965 1373 12142 1397
rect 12255 1444 12427 1533
rect -965 1293 12142 1317
rect -965 1241 2189 1293
rect 2241 1241 8697 1293
rect 8749 1241 12142 1293
rect -965 1217 12142 1241
rect -969 799 -813 811
rect -969 747 -945 799
rect -893 747 -813 799
rect -969 735 -813 747
rect 2121 799 2253 811
rect 2121 747 2189 799
rect 2241 747 2253 799
rect 2121 735 2253 747
rect 2309 799 2441 811
rect 2309 747 2321 799
rect 2373 747 2441 799
rect 2309 735 2441 747
rect 5375 735 5507 811
rect 5563 799 5695 811
rect 5563 747 5575 799
rect 5627 747 5695 799
rect 5563 735 5695 747
rect 8629 799 8761 811
rect 8629 747 8697 799
rect 8749 747 8761 799
rect 8629 735 8761 747
rect 8817 799 8949 811
rect 8817 747 8829 799
rect 8881 747 8949 799
rect 8817 735 8949 747
rect 11883 799 12195 811
rect 11883 747 12119 799
rect 12171 747 12195 799
rect 11883 735 12195 747
rect 2177 679 2253 735
tri 2253 679 2285 711 sw
rect 5431 679 5507 735
tri 5507 679 5539 711 sw
rect 8685 679 8761 735
tri 8761 679 8793 711 sw
tri 2177 571 2285 679 ne
tri 2285 579 2385 679 sw
rect 2285 571 2385 579
tri 5431 571 5539 679 ne
tri 5539 579 5639 679 sw
rect 5539 571 5639 579
tri 8685 571 8793 679 ne
tri 8793 579 8893 679 sw
rect 8793 571 8893 579
tri 2285 547 2309 571 ne
rect 2309 523 2385 571
tri 5539 547 5563 571 ne
rect 5563 523 5639 571
tri 8793 547 8817 571 ne
rect 8817 523 8893 571
rect -1125 511 -813 523
rect -1125 459 -1101 511
rect -1049 459 -813 511
rect -1125 447 -813 459
rect 2121 511 2253 523
rect 2121 459 2189 511
rect 2241 459 2253 511
rect 2121 447 2253 459
rect 2309 511 2441 523
rect 2309 459 2321 511
rect 2373 459 2441 511
rect 2309 447 2441 459
rect 5375 511 5507 523
rect 5375 459 5443 511
rect 5495 459 5507 511
rect 5375 447 5507 459
rect 5563 511 5695 523
rect 5563 459 5575 511
rect 5627 459 5695 511
rect 5563 447 5695 459
rect 8629 511 8761 523
rect 8629 459 8697 511
rect 8749 459 8761 511
rect 8629 447 8761 459
rect 8817 511 8949 523
rect 8817 459 8829 511
rect 8881 459 8949 511
rect 8817 447 8949 459
rect 11883 511 12039 523
rect 11883 459 11963 511
rect 12015 459 12039 511
rect 11883 447 12039 459
rect 2177 391 2253 447
tri 2253 391 2285 423 sw
rect 5431 391 5507 447
tri 5507 391 5539 423 sw
rect 8685 391 8761 447
tri 8761 391 8793 423 sw
tri 2177 283 2285 391 ne
tri 2285 291 2385 391 sw
rect 2285 283 2385 291
tri 5431 283 5539 391 ne
tri 5539 291 5639 391 sw
rect 5539 283 5639 291
tri 8685 283 8793 391 ne
tri 8793 291 8893 391 sw
rect 8793 283 8893 291
tri 2285 259 2309 283 ne
rect 2309 235 2385 283
tri 5539 259 5563 283 ne
rect 5563 235 5639 283
tri 8793 259 8817 283 ne
rect 8817 235 8893 283
rect -969 223 -813 235
rect -969 171 -945 223
rect -893 171 -813 223
rect -969 159 -813 171
rect 2121 223 2253 235
rect 2121 171 2189 223
rect 2241 171 2253 223
rect 2121 159 2253 171
rect 2309 223 2441 235
rect 2309 171 2321 223
rect 2373 171 2441 223
rect 2309 159 2441 171
rect 5375 223 5507 235
rect 5375 171 5443 223
rect 5495 171 5507 223
rect 5375 159 5507 171
rect 5563 223 5695 235
rect 5563 171 5575 223
rect 5627 171 5695 223
rect 5563 159 5695 171
rect 8629 223 8761 235
rect 8629 171 8697 223
rect 8749 171 8761 223
rect 8629 159 8761 171
rect 8817 223 8949 235
rect 8817 171 8829 223
rect 8881 171 8949 223
rect 8817 159 8949 171
rect 11883 223 12195 235
rect 11883 171 12119 223
rect 12171 171 12195 223
rect 11883 159 12195 171
rect 2177 103 2253 159
tri 2253 103 2285 135 sw
rect 5431 103 5507 159
tri 5507 103 5539 135 sw
rect 8685 103 8761 159
tri 8761 103 8793 135 sw
tri 2177 -5 2285 103 ne
tri 2285 3 2385 103 sw
rect 2285 -5 2385 3
tri 5431 -5 5539 103 ne
tri 5539 3 5639 103 sw
rect 5539 -5 5639 3
tri 8685 -5 8793 103 ne
tri 8793 3 8893 103 sw
rect 8793 -5 8893 3
tri 2285 -29 2309 -5 ne
rect 2309 -53 2385 -5
tri 5539 -29 5563 -5 ne
rect 5563 -53 5639 -5
tri 8793 -29 8817 -5 ne
rect 8817 -53 8893 -5
rect -1125 -65 -813 -53
rect -1125 -117 -1101 -65
rect -1049 -117 -813 -65
rect -1125 -129 -813 -117
rect 2121 -65 2253 -53
rect 2121 -117 2189 -65
rect 2241 -117 2253 -65
rect 2121 -129 2253 -117
rect 2309 -65 2441 -53
rect 2309 -117 2321 -65
rect 2373 -117 2441 -65
rect 2309 -129 2441 -117
rect 5375 -65 5507 -53
rect 5375 -117 5443 -65
rect 5495 -117 5507 -65
rect 5375 -129 5507 -117
rect 5563 -65 5695 -53
rect 5563 -117 5575 -65
rect 5627 -117 5695 -65
rect 5563 -129 5695 -117
rect 8629 -65 8761 -53
rect 8629 -117 8697 -65
rect 8749 -117 8761 -65
rect 8629 -129 8761 -117
rect 8817 -65 8949 -53
rect 8817 -117 8829 -65
rect 8881 -117 8949 -65
rect 8817 -129 8949 -117
rect 11883 -65 12039 -53
rect 11883 -117 11963 -65
rect 12015 -117 12039 -65
rect 11883 -129 12039 -117
rect 2177 -185 2253 -129
tri 2253 -185 2285 -153 sw
rect 5431 -185 5507 -129
tri 5507 -185 5539 -153 sw
rect 8685 -185 8761 -129
tri 8761 -185 8793 -153 sw
tri 2177 -293 2285 -185 ne
tri 2285 -285 2385 -185 sw
rect 2285 -293 2385 -285
tri 5431 -293 5539 -185 ne
tri 5539 -285 5639 -185 sw
rect 5539 -293 5639 -285
tri 8685 -293 8793 -185 ne
tri 8793 -285 8893 -185 sw
rect 8793 -293 8893 -285
tri 2285 -317 2309 -293 ne
rect 2309 -341 2385 -293
tri 5539 -317 5563 -293 ne
rect 5563 -341 5639 -293
tri 8793 -317 8817 -293 ne
rect 8817 -341 8893 -293
rect -969 -353 -813 -341
rect -969 -405 -945 -353
rect -893 -405 -813 -353
rect -969 -417 -813 -405
rect 2121 -353 2253 -341
rect 2121 -405 2189 -353
rect 2241 -405 2253 -353
rect 2121 -417 2253 -405
rect 2309 -417 2441 -341
rect 5375 -353 5507 -341
rect 5375 -405 5443 -353
rect 5495 -405 5507 -353
rect 5375 -417 5507 -405
rect 5563 -353 5695 -341
rect 5563 -405 5575 -353
rect 5627 -405 5695 -353
rect 5563 -417 5695 -405
rect 8629 -353 8761 -341
rect 8629 -405 8697 -353
rect 8749 -405 8761 -353
rect 8629 -417 8761 -405
rect 8817 -417 8949 -341
rect 11883 -353 12195 -341
rect 11883 -405 12119 -353
rect 12171 -405 12195 -353
rect 11883 -417 12195 -405
rect -1125 -847 12195 -823
rect -1125 -899 -1101 -847
rect -1049 -899 5443 -847
rect 5495 -899 12119 -847
rect 12171 -899 12195 -847
rect -1125 -923 12195 -899
rect -1357 -1139 -1185 -1050
rect -969 -1003 12039 -979
rect -969 -1055 -946 -1003
rect -894 -1055 5575 -1003
rect 5627 -1055 11964 -1003
rect 12016 -1055 12039 -1003
rect -969 -1079 12039 -1055
rect 12255 -1050 12318 1444
rect 12364 -1050 12427 1444
rect 12255 -1139 12427 -1050
rect -1357 -1199 12427 -1139
rect -1357 -1202 -801 -1199
rect -749 -1202 2057 -1199
rect 2109 -1202 2453 -1199
rect 2505 -1202 5311 -1199
rect 5363 -1202 5707 -1199
rect 5759 -1202 8565 -1199
rect 8617 -1202 8961 -1199
rect 9013 -1202 11819 -1199
rect 11871 -1202 12427 -1199
rect -1357 -1248 -1169 -1202
rect 12239 -1248 12427 -1202
rect -1357 -1251 -801 -1248
rect -749 -1251 2057 -1248
rect 2109 -1251 2453 -1248
rect 2505 -1251 5311 -1248
rect 5363 -1251 5707 -1248
rect 5759 -1251 8565 -1248
rect 8617 -1251 8961 -1248
rect 9013 -1251 11819 -1248
rect 11871 -1251 12427 -1248
rect -1357 -1311 12427 -1251
<< via1 >>
rect -801 1642 -749 1645
rect 2057 1642 2109 1645
rect 2453 1642 2505 1645
rect 5311 1642 5363 1645
rect 5707 1642 5759 1645
rect 8565 1642 8617 1645
rect 8961 1642 9013 1645
rect 11819 1642 11871 1645
rect -801 1596 -749 1642
rect 2057 1596 2109 1642
rect 2453 1596 2505 1642
rect 5311 1596 5363 1642
rect 5707 1596 5759 1642
rect 8565 1596 8617 1642
rect 8961 1596 9013 1642
rect 11819 1596 11871 1642
rect -801 1593 -749 1596
rect 2057 1593 2109 1596
rect 2453 1593 2505 1596
rect 5311 1593 5363 1596
rect 5707 1593 5759 1596
rect 8565 1593 8617 1596
rect 8961 1593 9013 1596
rect 11819 1593 11871 1596
rect 2321 1397 2373 1449
rect 8829 1397 8881 1449
rect 2189 1241 2241 1293
rect 8697 1241 8749 1293
rect -801 1035 -749 1087
rect 2057 1035 2109 1087
rect 2453 1035 2505 1087
rect 5311 1035 5363 1087
rect 5707 1035 5759 1087
rect 8565 1035 8617 1087
rect 8961 1035 9013 1087
rect 11819 1035 11871 1087
rect -945 747 -893 799
rect 2189 747 2241 799
rect 2321 747 2373 799
rect 5575 747 5627 799
rect 8697 747 8749 799
rect 8829 747 8881 799
rect 12119 747 12171 799
rect -1101 459 -1049 511
rect 2189 459 2241 511
rect 2321 459 2373 511
rect 5443 459 5495 511
rect 5575 459 5627 511
rect 8697 459 8749 511
rect 8829 459 8881 511
rect 11963 459 12015 511
rect -945 171 -893 223
rect 2189 171 2241 223
rect 2321 171 2373 223
rect 5443 171 5495 223
rect 5575 171 5627 223
rect 8697 171 8749 223
rect 8829 171 8881 223
rect 12119 171 12171 223
rect -1101 -117 -1049 -65
rect 2189 -117 2241 -65
rect 2321 -117 2373 -65
rect 5443 -117 5495 -65
rect 5575 -117 5627 -65
rect 8697 -117 8749 -65
rect 8829 -117 8881 -65
rect 11963 -117 12015 -65
rect -945 -405 -893 -353
rect 2189 -405 2241 -353
rect 5443 -405 5495 -353
rect 5575 -405 5627 -353
rect 8697 -405 8749 -353
rect 12119 -405 12171 -353
rect -801 -693 -749 -641
rect 2057 -693 2109 -641
rect 2453 -693 2505 -641
rect 5311 -693 5363 -641
rect 5707 -693 5759 -641
rect 8565 -693 8617 -641
rect 8961 -693 9013 -641
rect 11819 -693 11871 -641
rect -1101 -899 -1049 -847
rect 5443 -899 5495 -847
rect 12119 -899 12171 -847
rect -946 -1055 -894 -1003
rect 5575 -1055 5627 -1003
rect 11964 -1055 12016 -1003
rect -801 -1202 -749 -1199
rect 2057 -1202 2109 -1199
rect 2453 -1202 2505 -1199
rect 5311 -1202 5363 -1199
rect 5707 -1202 5759 -1199
rect 8565 -1202 8617 -1199
rect 8961 -1202 9013 -1199
rect 11819 -1202 11871 -1199
rect -801 -1248 -749 -1202
rect 2057 -1248 2109 -1202
rect 2453 -1248 2505 -1202
rect 5311 -1248 5363 -1202
rect 5707 -1248 5759 -1202
rect 8565 -1248 8617 -1202
rect 8961 -1248 9013 -1202
rect 11819 -1248 11871 -1202
rect -801 -1251 -749 -1248
rect 2057 -1251 2109 -1248
rect 2453 -1251 2505 -1248
rect 5311 -1251 5363 -1248
rect 5707 -1251 5759 -1248
rect 8565 -1251 8617 -1248
rect 8961 -1251 9013 -1248
rect 11819 -1251 11871 -1248
<< metal2 >>
rect -813 1645 -737 1647
rect -813 1593 -801 1645
rect -749 1593 -737 1645
rect -813 1087 -737 1593
rect -813 1035 -801 1087
rect -749 1035 -737 1087
rect -813 1023 -737 1035
rect 2045 1645 2121 1647
rect 2045 1593 2057 1645
rect 2109 1593 2121 1645
rect 2045 1087 2121 1593
rect 2441 1645 2517 1647
rect 2441 1593 2453 1645
rect 2505 1593 2517 1645
rect 2309 1449 2385 1473
rect 2309 1397 2321 1449
rect 2373 1397 2385 1449
rect 2045 1035 2057 1087
rect 2109 1035 2121 1087
rect 2045 1023 2121 1035
rect 2177 1293 2253 1317
rect 2177 1241 2189 1293
rect 2241 1241 2253 1293
rect -969 799 -869 811
rect -969 747 -945 799
rect -893 747 -869 799
rect -1125 511 -1025 523
rect -1125 459 -1101 511
rect -1049 459 -1025 511
rect -1125 -65 -1025 459
rect -1125 -117 -1101 -65
rect -1049 -117 -1025 -65
rect -1125 -847 -1025 -117
rect -1125 -899 -1101 -847
rect -1049 -899 -1025 -847
rect -1125 -923 -1025 -899
rect -969 223 -869 747
rect 2177 799 2253 1241
rect 2177 747 2189 799
rect 2241 747 2253 799
rect 2177 735 2253 747
rect 2309 799 2385 1397
rect 2441 1087 2517 1593
rect 2441 1035 2453 1087
rect 2505 1035 2517 1087
rect 2441 1023 2517 1035
rect 5299 1645 5375 1647
rect 5299 1593 5311 1645
rect 5363 1593 5375 1645
rect 5299 1087 5375 1593
rect 5299 1035 5311 1087
rect 5363 1035 5375 1087
rect 5299 1023 5375 1035
rect 5695 1645 5771 1647
rect 5695 1593 5707 1645
rect 5759 1593 5771 1645
rect 5695 1087 5771 1593
rect 5695 1035 5707 1087
rect 5759 1035 5771 1087
rect 5695 1023 5771 1035
rect 8553 1645 8629 1647
rect 8553 1593 8565 1645
rect 8617 1593 8629 1645
rect 8553 1087 8629 1593
rect 8949 1645 9025 1647
rect 8949 1593 8961 1645
rect 9013 1593 9025 1645
rect 8817 1449 8893 1473
rect 8817 1397 8829 1449
rect 8881 1397 8893 1449
rect 8553 1035 8565 1087
rect 8617 1035 8629 1087
rect 8553 1023 8629 1035
rect 8685 1293 8761 1317
rect 8685 1241 8697 1293
rect 8749 1241 8761 1293
rect 2309 747 2321 799
rect 2373 747 2385 799
tri 2201 603 2309 711 se
rect 2309 679 2385 747
rect 5563 799 5639 811
rect 5563 747 5575 799
rect 5627 747 5639 799
tri 2309 603 2385 679 nw
tri 5455 603 5563 711 se
rect 5563 679 5639 747
rect 8685 799 8761 1241
rect 8685 747 8697 799
rect 8749 747 8761 799
rect 8685 735 8761 747
rect 8817 799 8893 1397
rect 8949 1087 9025 1593
rect 8949 1035 8961 1087
rect 9013 1035 9025 1087
rect 8949 1023 9025 1035
rect 11807 1645 11883 1647
rect 11807 1593 11819 1645
rect 11871 1593 11883 1645
rect 11807 1087 11883 1593
rect 11807 1035 11819 1087
rect 11871 1035 11883 1087
rect 11807 1023 11883 1035
rect 8817 747 8829 799
rect 8881 747 8893 799
tri 5563 603 5639 679 nw
tri 8709 603 8817 711 se
rect 8817 679 8893 747
tri 8817 603 8893 679 nw
rect 12095 799 12195 811
rect 12095 747 12119 799
rect 12171 747 12195 799
tri 2177 579 2201 603 se
rect 2201 579 2253 603
rect 2177 511 2253 579
tri 2253 547 2309 603 nw
tri 5431 579 5455 603 se
rect 5455 579 5507 603
rect 2177 459 2189 511
rect 2241 459 2253 511
rect 2177 447 2253 459
rect 2309 511 2385 523
rect 2309 459 2321 511
rect 2373 459 2385 511
tri 2201 315 2309 423 se
rect 2309 391 2385 459
rect 5431 511 5507 579
tri 5507 547 5563 603 nw
tri 8685 579 8709 603 se
rect 8709 579 8761 603
rect 5431 459 5443 511
rect 5495 459 5507 511
rect 5431 447 5507 459
rect 5563 511 5639 523
rect 5563 459 5575 511
rect 5627 459 5639 511
tri 2309 315 2385 391 nw
tri 5455 315 5563 423 se
rect 5563 391 5639 459
rect 8685 511 8761 579
tri 8761 547 8817 603 nw
rect 8685 459 8697 511
rect 8749 459 8761 511
rect 8685 447 8761 459
rect 8817 511 8893 523
rect 8817 459 8829 511
rect 8881 459 8893 511
tri 5563 315 5639 391 nw
tri 8709 315 8817 423 se
rect 8817 391 8893 459
tri 8817 315 8893 391 nw
rect 11939 511 12039 523
rect 11939 459 11963 511
rect 12015 459 12039 511
rect -969 171 -945 223
rect -893 171 -869 223
rect -969 -353 -869 171
tri 2177 291 2201 315 se
rect 2201 291 2253 315
rect 2177 223 2253 291
tri 2253 259 2309 315 nw
tri 5431 291 5455 315 se
rect 5455 291 5507 315
rect 2177 171 2189 223
rect 2241 171 2253 223
rect 2177 159 2253 171
rect 2309 223 2385 235
rect 2309 171 2321 223
rect 2373 171 2385 223
tri 2201 27 2309 135 se
rect 2309 103 2385 171
rect 5431 223 5507 291
tri 5507 259 5563 315 nw
tri 8685 291 8709 315 se
rect 8709 291 8761 315
rect 5431 171 5443 223
rect 5495 171 5507 223
rect 5431 159 5507 171
rect 5563 223 5639 235
rect 5563 171 5575 223
rect 5627 171 5639 223
tri 2309 27 2385 103 nw
tri 5455 27 5563 135 se
rect 5563 103 5639 171
rect 8685 223 8761 291
tri 8761 259 8817 315 nw
rect 8685 171 8697 223
rect 8749 171 8761 223
rect 8685 159 8761 171
rect 8817 223 8893 235
rect 8817 171 8829 223
rect 8881 171 8893 223
tri 5563 27 5639 103 nw
tri 8709 27 8817 135 se
rect 8817 103 8893 171
tri 8817 27 8893 103 nw
tri 2177 3 2201 27 se
rect 2201 3 2253 27
rect 2177 -65 2253 3
tri 2253 -29 2309 27 nw
tri 5431 3 5455 27 se
rect 5455 3 5507 27
rect 2177 -117 2189 -65
rect 2241 -117 2253 -65
rect 2177 -129 2253 -117
rect 2309 -65 2385 -53
rect 2309 -117 2321 -65
rect 2373 -117 2385 -65
tri 2201 -261 2309 -153 se
rect 2309 -185 2385 -117
rect 5431 -65 5507 3
tri 5507 -29 5563 27 nw
tri 8685 3 8709 27 se
rect 8709 3 8761 27
rect 5431 -117 5443 -65
rect 5495 -117 5507 -65
rect 5431 -129 5507 -117
rect 5563 -65 5639 -53
rect 5563 -117 5575 -65
rect 5627 -117 5639 -65
tri 2309 -261 2385 -185 nw
tri 5455 -261 5563 -153 se
rect 5563 -185 5639 -117
rect 8685 -65 8761 3
tri 8761 -29 8817 27 nw
rect 8685 -117 8697 -65
rect 8749 -117 8761 -65
rect 8685 -129 8761 -117
rect 8817 -65 8893 -53
rect 8817 -117 8829 -65
rect 8881 -117 8893 -65
tri 5563 -261 5639 -185 nw
tri 8709 -261 8817 -153 se
rect 8817 -185 8893 -117
tri 8817 -261 8893 -185 nw
rect 11939 -65 12039 459
rect 11939 -117 11963 -65
rect 12015 -117 12039 -65
rect -969 -405 -945 -353
rect -893 -405 -869 -353
rect -969 -1003 -869 -405
tri 2177 -285 2201 -261 se
rect 2201 -285 2253 -261
rect 2177 -353 2253 -285
tri 2253 -317 2309 -261 nw
tri 5431 -285 5455 -261 se
rect 5455 -285 5507 -261
rect 2177 -405 2189 -353
rect 2241 -405 2253 -353
rect 2177 -417 2253 -405
rect 5431 -353 5507 -285
tri 5507 -317 5563 -261 nw
tri 8685 -285 8709 -261 se
rect 8709 -285 8761 -261
rect 5431 -405 5443 -353
rect 5495 -405 5507 -353
rect -969 -1055 -946 -1003
rect -894 -1055 -869 -1003
rect -969 -1079 -869 -1055
rect -813 -641 -737 -629
rect -813 -693 -801 -641
rect -749 -693 -737 -641
rect -813 -1199 -737 -693
rect -813 -1251 -801 -1199
rect -749 -1251 -737 -1199
rect -813 -1253 -737 -1251
rect 2045 -641 2121 -629
rect 2045 -693 2057 -641
rect 2109 -693 2121 -641
rect 2045 -1199 2121 -693
rect 2045 -1251 2057 -1199
rect 2109 -1251 2121 -1199
rect 2045 -1253 2121 -1251
rect 2441 -641 2517 -629
rect 2441 -693 2453 -641
rect 2505 -693 2517 -641
rect 2441 -1199 2517 -693
rect 2441 -1251 2453 -1199
rect 2505 -1251 2517 -1199
rect 2441 -1253 2517 -1251
rect 5299 -641 5375 -629
rect 5299 -693 5311 -641
rect 5363 -693 5375 -641
rect 5299 -1199 5375 -693
rect 5431 -847 5507 -405
rect 5431 -899 5443 -847
rect 5495 -899 5507 -847
rect 5431 -923 5507 -899
rect 5563 -353 5639 -341
rect 5563 -405 5575 -353
rect 5627 -405 5639 -353
rect 5563 -1003 5639 -405
rect 8685 -353 8761 -285
tri 8761 -317 8817 -261 nw
rect 8685 -405 8697 -353
rect 8749 -405 8761 -353
rect 8685 -417 8761 -405
rect 5563 -1055 5575 -1003
rect 5627 -1055 5639 -1003
rect 5563 -1079 5639 -1055
rect 5695 -641 5771 -629
rect 5695 -693 5707 -641
rect 5759 -693 5771 -641
rect 5299 -1251 5311 -1199
rect 5363 -1251 5375 -1199
rect 5299 -1253 5375 -1251
rect 5695 -1199 5771 -693
rect 5695 -1251 5707 -1199
rect 5759 -1251 5771 -1199
rect 5695 -1253 5771 -1251
rect 8553 -641 8629 -629
rect 8553 -693 8565 -641
rect 8617 -693 8629 -641
rect 8553 -1199 8629 -693
rect 8553 -1251 8565 -1199
rect 8617 -1251 8629 -1199
rect 8553 -1253 8629 -1251
rect 8949 -641 9025 -629
rect 8949 -693 8961 -641
rect 9013 -693 9025 -641
rect 8949 -1199 9025 -693
rect 8949 -1251 8961 -1199
rect 9013 -1251 9025 -1199
rect 8949 -1253 9025 -1251
rect 11807 -641 11883 -629
rect 11807 -693 11819 -641
rect 11871 -693 11883 -641
rect 11807 -1199 11883 -693
rect 11939 -1003 12039 -117
rect 12095 223 12195 747
rect 12095 171 12119 223
rect 12171 171 12195 223
rect 12095 -353 12195 171
rect 12095 -405 12119 -353
rect 12171 -405 12195 -353
rect 12095 -847 12195 -405
rect 12095 -899 12119 -847
rect 12171 -899 12195 -847
rect 12095 -923 12195 -899
rect 11939 -1055 11964 -1003
rect 12016 -1055 12039 -1003
rect 11939 -1079 12039 -1055
rect 11807 -1251 11819 -1199
rect 11871 -1251 11883 -1199
rect 11807 -1253 11883 -1251
use res_13p37u  res_13p37u_0
timestamp 1586907467
transform 1 0 8871 0 1 881
box 78 80 3012 280
use res_13p37u  res_13p37u_1
timestamp 1586907467
transform 1 0 8871 0 1 593
box 78 80 3012 280
use res_13p37u  res_13p37u_2
timestamp 1586907467
transform 1 0 8871 0 1 305
box 78 80 3012 280
use res_13p37u  res_13p37u_3
timestamp 1586907467
transform 1 0 8871 0 1 17
box 78 80 3012 280
use res_13p37u  res_13p37u_4
timestamp 1586907467
transform 1 0 8871 0 1 -271
box 78 80 3012 280
use res_13p37u  res_13p37u_5
timestamp 1586907467
transform 1 0 8871 0 1 -559
box 78 80 3012 280
use res_13p37u  res_13p37u_6
timestamp 1586907467
transform 1 0 8871 0 1 -847
box 78 80 3012 280
use res_13p37u  res_13p37u_7
timestamp 1586907467
transform 1 0 5617 0 1 881
box 78 80 3012 280
use res_13p37u  res_13p37u_8
timestamp 1586907467
transform 1 0 5617 0 1 593
box 78 80 3012 280
use res_13p37u  res_13p37u_9
timestamp 1586907467
transform 1 0 5617 0 1 305
box 78 80 3012 280
use res_13p37u  res_13p37u_10
timestamp 1586907467
transform 1 0 5617 0 1 17
box 78 80 3012 280
use res_13p37u  res_13p37u_11
timestamp 1586907467
transform 1 0 5617 0 1 -271
box 78 80 3012 280
use res_13p37u  res_13p37u_12
timestamp 1586907467
transform 1 0 5617 0 1 -559
box 78 80 3012 280
use res_13p37u  res_13p37u_13
timestamp 1586907467
transform 1 0 5617 0 1 -847
box 78 80 3012 280
use res_13p37u  res_13p37u_14
timestamp 1586907467
transform 1 0 2363 0 1 -847
box 78 80 3012 280
use res_13p37u  res_13p37u_15
timestamp 1586907467
transform 1 0 -891 0 1 -847
box 78 80 3012 280
use res_13p37u  res_13p37u_16
timestamp 1586907467
transform 1 0 2363 0 1 -559
box 78 80 3012 280
use res_13p37u  res_13p37u_17
timestamp 1586907467
transform 1 0 -891 0 1 -559
box 78 80 3012 280
use res_13p37u  res_13p37u_18
timestamp 1586907467
transform 1 0 -891 0 1 17
box 78 80 3012 280
use res_13p37u  res_13p37u_19
timestamp 1586907467
transform 1 0 2363 0 1 -271
box 78 80 3012 280
use res_13p37u  res_13p37u_20
timestamp 1586907467
transform 1 0 -891 0 1 -271
box 78 80 3012 280
use res_13p37u  res_13p37u_21
timestamp 1586907467
transform 1 0 2363 0 1 17
box 78 80 3012 280
use res_13p37u  res_13p37u_22
timestamp 1586907467
transform 1 0 -891 0 1 305
box 78 80 3012 280
use res_13p37u  res_13p37u_23
timestamp 1586907467
transform 1 0 2363 0 1 305
box 78 80 3012 280
use res_13p37u  res_13p37u_24
timestamp 1586907467
transform 1 0 2363 0 1 593
box 78 80 3012 280
use res_13p37u  res_13p37u_25
timestamp 1586907467
transform 1 0 -891 0 1 593
box 78 80 3012 280
use res_13p37u  res_13p37u_26
timestamp 1586907467
transform 1 0 2363 0 1 881
box 78 80 3012 280
use res_13p37u  res_13p37u_27
timestamp 1586907467
transform 1 0 -891 0 1 881
box 78 80 3012 280
<< labels >>
flabel metal1 s -1284 1591 -1284 1591 2 FreeSans 600 0 0 0 VSS
port 1 nsew
flabel metal1 s -945 1254 -945 1254 2 FreeSans 600 0 0 0 A1
port 2 nsew
flabel metal1 s -951 1394 -951 1394 2 FreeSans 600 0 0 0 A2
port 3 nsew
flabel metal1 s -849 -911 -849 -911 2 FreeSans 600 0 0 0 B2
port 4 nsew
flabel metal1 s -832 -1056 -832 -1056 2 FreeSans 600 0 0 0 B1
port 5 nsew
<< properties >>
string path 27.345 2.235 27.345 2.815 28.005 3.475 28.005 4.055 
<< end >>
