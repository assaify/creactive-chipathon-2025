magic
tech gf180mcuD
magscale 1 10
timestamp 1757676927
<< error_s >>
rect -1366 -1582 -1364 -1572
rect -1364 -1592 -1354 -1582
rect -1368 -1638 -1366 -1636
rect -1364 -1638 -1354 -1628
rect -1368 -1648 -1364 -1638
rect -1368 -1777 -1366 -1648
rect 990 -1697 1101 -936
rect -756 -1884 -754 -1740
rect -758 -1894 -754 -1884
rect -768 -1904 -758 -1894
rect -756 -1896 -754 -1894
rect -768 -1950 -758 -1940
rect -758 -1960 -756 -1950
rect -1368 -3069 -1366 -2938
rect 415 -3294 417 -3016
rect 2170 -3292 2172 -3032
<< metal1 >>
rect -1641 -864 4570 -664
rect -1450 -1052 -1250 -864
rect 895 -1232 1066 -1052
rect 1004 -2524 1119 -2344
rect -1641 -3374 4570 -3352
rect -1641 -3530 -1074 -3374
rect -918 -3530 4570 -3374
rect -1641 -3552 4570 -3530
<< via1 >>
rect -1074 -2228 -918 -2072
rect -1074 -3530 -918 -3374
<< metal2 >>
rect 916 -1893 1016 -1872
rect 916 -1949 938 -1893
rect 994 -1949 1016 -1893
rect -1096 -2072 -896 -2060
rect -1096 -2228 -1074 -2072
rect -918 -2228 -896 -2072
rect -1096 -3374 -896 -2228
rect 916 -2600 1016 -1949
rect 916 -2656 938 -2600
rect 994 -2656 1016 -2600
rect 916 -2678 1016 -2656
rect -1096 -3530 -1074 -3374
rect -918 -3530 -896 -3374
rect -1096 -3552 -896 -3530
<< via2 >>
rect 938 -1949 994 -1893
rect 938 -2656 994 -2600
<< metal3 >>
rect -1641 -1660 4570 -1560
rect -1641 -1816 4570 -1716
rect -1641 -1972 -569 -1872
rect 616 -1893 4570 -1872
rect 616 -1949 938 -1893
rect 994 -1949 4570 -1893
rect 616 -1972 4570 -1949
rect 916 -2600 1119 -2578
rect 916 -2656 938 -2600
rect 994 -2656 1119 -2600
rect 916 -2678 1119 -2656
rect -1641 -2834 4570 -2734
<< via3 >>
rect 1827 -1130 2195 -970
rect 1280 -1428 1648 -1268
<< metal4 >>
rect 1264 -1268 1664 -636
rect 1811 -918 2211 -850
rect 1811 -1182 1827 -918
rect 2195 -1182 2211 -918
rect 1811 -1250 2211 -1182
rect 1264 -1428 1280 -1268
rect 1648 -1428 1664 -1268
rect 1264 -3580 1664 -1428
<< via4 >>
rect 1827 -970 2195 -918
rect 1827 -1130 2195 -970
rect 1827 -1182 2195 -1130
<< metal5 >>
rect -1641 -918 4570 -850
rect -1641 -1182 1827 -918
rect 2195 -1182 4570 -918
rect -1641 -1250 4570 -1182
use dff_2ph_clk$1  dff_2ph_clk$1_0
timestamp 1757676927
transform 1 0 671 0 1 -1142
box -2326 -2405 310 103
use gf180mcu_fd_sc_mcu9t5v0__fill_2  gf180mcu_fd_sc_mcu9t5v0__fill_2_0
timestamp 1757676927
transform 1 0 895 0 1 -3442
box -86 -90 310 1098
use tgate$1  tgate$1_0
timestamp 1757676927
transform 1 0 2290 0 1 -2234
box -1300 -1318 2256 1570
<< labels >>
flabel metal1 s -1638 -3452 -1638 -3452 2 FreeSans 73 0 0 0 VSSD
port 1 nsew
flabel metal1 s -1638 -764 -1638 -764 2 FreeSans 73 0 0 0 VDDD
port 2 nsew
flabel metal3 s 2522 -1348 2522 -1348 2 FreeSans 89 0 0 0 T2
port 3 nsew
flabel metal3 s -1638 -2784 -1638 -2784 2 FreeSans 89 0 0 0 EN
port 4 nsew
flabel metal3 s 2522 -1050 2522 -1050 2 FreeSans 89 0 0 0 T1
port 5 nsew
flabel metal3 s -801 -1922 -801 -1922 2 FreeSans 89 0 0 0 DATA_IN
port 6 nsew
flabel metal3 s -801 -1766 -801 -1766 2 FreeSans 89 0 0 0 CLK_PH2
port 7 nsew
flabel metal3 s -801 -1610 -801 -1610 2 FreeSans 89 0 0 0 CLK_PH1
port 8 nsew
flabel metal3 s 4567 -1922 4567 -1922 8 FreeSans 89 0 0 0 DATA_OUT
port 9 nsew
<< properties >>
string path -8.205 -5.250 22.850 -5.250 
<< end >>
