magic
tech gf180mcuD
magscale 1 10
timestamp 1755276408
<< nwell >>
rect -350 -4558 350 4558
<< pmos >>
rect -100 2348 100 4348
rect -100 116 100 2116
rect -100 -2116 100 -116
rect -100 -4348 100 -2348
<< pdiff >>
rect -188 4335 -100 4348
rect -188 2361 -175 4335
rect -129 2361 -100 4335
rect -188 2348 -100 2361
rect 100 4335 188 4348
rect 100 2361 129 4335
rect 175 2361 188 4335
rect 100 2348 188 2361
rect -188 2103 -100 2116
rect -188 129 -175 2103
rect -129 129 -100 2103
rect -188 116 -100 129
rect 100 2103 188 2116
rect 100 129 129 2103
rect 175 129 188 2103
rect 100 116 188 129
rect -188 -129 -100 -116
rect -188 -2103 -175 -129
rect -129 -2103 -100 -129
rect -188 -2116 -100 -2103
rect 100 -129 188 -116
rect 100 -2103 129 -129
rect 175 -2103 188 -129
rect 100 -2116 188 -2103
rect -188 -2361 -100 -2348
rect -188 -4335 -175 -2361
rect -129 -4335 -100 -2361
rect -188 -4348 -100 -4335
rect 100 -2361 188 -2348
rect 100 -4335 129 -2361
rect 175 -4335 188 -2361
rect 100 -4348 188 -4335
<< pdiffc >>
rect -175 2361 -129 4335
rect 129 2361 175 4335
rect -175 129 -129 2103
rect 129 129 175 2103
rect -175 -2103 -129 -129
rect 129 -2103 175 -129
rect -175 -4335 -129 -2361
rect 129 -4335 175 -2361
<< nsubdiff >>
rect -326 4462 326 4534
rect -326 4418 -254 4462
rect -326 -4418 -313 4418
rect -267 -4418 -254 4418
rect 254 4418 326 4462
rect -326 -4462 -254 -4418
rect 254 -4418 267 4418
rect 313 -4418 326 4418
rect 254 -4462 326 -4418
rect -326 -4534 326 -4462
<< nsubdiffcont >>
rect -313 -4418 -267 4418
rect 267 -4418 313 4418
<< polysilicon >>
rect -100 4427 100 4440
rect -100 4381 -87 4427
rect 87 4381 100 4427
rect -100 4348 100 4381
rect -100 2315 100 2348
rect -100 2269 -87 2315
rect 87 2269 100 2315
rect -100 2256 100 2269
rect -100 2195 100 2208
rect -100 2149 -87 2195
rect 87 2149 100 2195
rect -100 2116 100 2149
rect -100 83 100 116
rect -100 37 -87 83
rect 87 37 100 83
rect -100 24 100 37
rect -100 -37 100 -24
rect -100 -83 -87 -37
rect 87 -83 100 -37
rect -100 -116 100 -83
rect -100 -2149 100 -2116
rect -100 -2195 -87 -2149
rect 87 -2195 100 -2149
rect -100 -2208 100 -2195
rect -100 -2269 100 -2256
rect -100 -2315 -87 -2269
rect 87 -2315 100 -2269
rect -100 -2348 100 -2315
rect -100 -4381 100 -4348
rect -100 -4427 -87 -4381
rect 87 -4427 100 -4381
rect -100 -4440 100 -4427
<< polycontact >>
rect -87 4381 87 4427
rect -87 2269 87 2315
rect -87 2149 87 2195
rect -87 37 87 83
rect -87 -83 87 -37
rect -87 -2195 87 -2149
rect -87 -2315 87 -2269
rect -87 -4427 87 -4381
<< metal1 >>
rect -313 4475 313 4521
rect -313 4418 -267 4475
rect -98 4381 -87 4427
rect 87 4381 98 4427
rect 267 4418 313 4475
rect -175 4335 -129 4346
rect -175 2350 -129 2361
rect 129 4335 175 4346
rect 129 2350 175 2361
rect -98 2269 -87 2315
rect 87 2269 98 2315
rect -98 2149 -87 2195
rect 87 2149 98 2195
rect -175 2103 -129 2114
rect -175 118 -129 129
rect 129 2103 175 2114
rect 129 118 175 129
rect -98 37 -87 83
rect 87 37 98 83
rect -98 -83 -87 -37
rect 87 -83 98 -37
rect -175 -129 -129 -118
rect -175 -2114 -129 -2103
rect 129 -129 175 -118
rect 129 -2114 175 -2103
rect -98 -2195 -87 -2149
rect 87 -2195 98 -2149
rect -98 -2315 -87 -2269
rect 87 -2315 98 -2269
rect -175 -2361 -129 -2350
rect -175 -4346 -129 -4335
rect 129 -2361 175 -2350
rect 129 -4346 175 -4335
rect -313 -4475 -267 -4418
rect -98 -4427 -87 -4381
rect 87 -4427 98 -4381
rect 267 -4475 313 -4418
rect -313 -4521 313 -4475
<< properties >>
string FIXED_BBOX -290 -4498 290 4498
string gencell pfet_03v3
string library gf180mcu
string parameters w 10.0 l 1.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 class mosfet full_metal 1 compatible {pfet_03v3 pfet_06v0} ad {int((nf+1)/2) * W/nf * 0.18u} as {int((nf+2)/2) * W/nf * 0.18u} pd {2*int((nf+1)/2) * (W/nf + 0.18u)} ps {2*int((nf+2)/2) * (W/nf + 0.18u)} nrd {0.18u / W} nrs {0.18u / W} sa 0 sb 0 sd 0
<< end >>
