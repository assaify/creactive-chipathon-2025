magic
tech gf180mcuD
magscale 1 10
timestamp 1755280221
<< mimcap >>
rect -17567 7900 -16567 7980
rect -17567 7060 -17487 7900
rect -16647 7060 -16567 7900
rect -17567 6980 -16567 7060
rect -15953 7900 -14953 7980
rect -15953 7060 -15873 7900
rect -15033 7060 -14953 7900
rect -15953 6980 -14953 7060
rect -14339 7900 -13339 7980
rect -14339 7060 -14259 7900
rect -13419 7060 -13339 7900
rect -14339 6980 -13339 7060
rect -12725 7900 -11725 7980
rect -12725 7060 -12645 7900
rect -11805 7060 -11725 7900
rect -12725 6980 -11725 7060
rect -11111 7900 -10111 7980
rect -11111 7060 -11031 7900
rect -10191 7060 -10111 7900
rect -11111 6980 -10111 7060
rect -9497 7900 -8497 7980
rect -9497 7060 -9417 7900
rect -8577 7060 -8497 7900
rect -9497 6980 -8497 7060
rect -7883 7900 -6883 7980
rect -7883 7060 -7803 7900
rect -6963 7060 -6883 7900
rect -7883 6980 -6883 7060
rect -6269 7900 -5269 7980
rect -6269 7060 -6189 7900
rect -5349 7060 -5269 7900
rect -6269 6980 -5269 7060
rect -4655 7900 -3655 7980
rect -4655 7060 -4575 7900
rect -3735 7060 -3655 7900
rect -4655 6980 -3655 7060
rect -3041 7900 -2041 7980
rect -3041 7060 -2961 7900
rect -2121 7060 -2041 7900
rect -3041 6980 -2041 7060
rect -1427 7900 -427 7980
rect -1427 7060 -1347 7900
rect -507 7060 -427 7900
rect -1427 6980 -427 7060
rect 187 7900 1187 7980
rect 187 7060 267 7900
rect 1107 7060 1187 7900
rect 187 6980 1187 7060
rect 1801 7900 2801 7980
rect 1801 7060 1881 7900
rect 2721 7060 2801 7900
rect 1801 6980 2801 7060
rect 3415 7900 4415 7980
rect 3415 7060 3495 7900
rect 4335 7060 4415 7900
rect 3415 6980 4415 7060
rect 5029 7900 6029 7980
rect 5029 7060 5109 7900
rect 5949 7060 6029 7900
rect 5029 6980 6029 7060
rect 6643 7900 7643 7980
rect 6643 7060 6723 7900
rect 7563 7060 7643 7900
rect 6643 6980 7643 7060
rect 8257 7900 9257 7980
rect 8257 7060 8337 7900
rect 9177 7060 9257 7900
rect 8257 6980 9257 7060
rect 9871 7900 10871 7980
rect 9871 7060 9951 7900
rect 10791 7060 10871 7900
rect 9871 6980 10871 7060
rect 11485 7900 12485 7980
rect 11485 7060 11565 7900
rect 12405 7060 12485 7900
rect 11485 6980 12485 7060
rect 13099 7900 14099 7980
rect 13099 7060 13179 7900
rect 14019 7060 14099 7900
rect 13099 6980 14099 7060
rect 14713 7900 15713 7980
rect 14713 7060 14793 7900
rect 15633 7060 15713 7900
rect 14713 6980 15713 7060
rect 16327 7900 17327 7980
rect 16327 7060 16407 7900
rect 17247 7060 17327 7900
rect 16327 6980 17327 7060
rect -17567 6540 -16567 6620
rect -17567 5700 -17487 6540
rect -16647 5700 -16567 6540
rect -17567 5620 -16567 5700
rect -15953 6540 -14953 6620
rect -15953 5700 -15873 6540
rect -15033 5700 -14953 6540
rect -15953 5620 -14953 5700
rect -14339 6540 -13339 6620
rect -14339 5700 -14259 6540
rect -13419 5700 -13339 6540
rect -14339 5620 -13339 5700
rect -12725 6540 -11725 6620
rect -12725 5700 -12645 6540
rect -11805 5700 -11725 6540
rect -12725 5620 -11725 5700
rect -11111 6540 -10111 6620
rect -11111 5700 -11031 6540
rect -10191 5700 -10111 6540
rect -11111 5620 -10111 5700
rect -9497 6540 -8497 6620
rect -9497 5700 -9417 6540
rect -8577 5700 -8497 6540
rect -9497 5620 -8497 5700
rect -7883 6540 -6883 6620
rect -7883 5700 -7803 6540
rect -6963 5700 -6883 6540
rect -7883 5620 -6883 5700
rect -6269 6540 -5269 6620
rect -6269 5700 -6189 6540
rect -5349 5700 -5269 6540
rect -6269 5620 -5269 5700
rect -4655 6540 -3655 6620
rect -4655 5700 -4575 6540
rect -3735 5700 -3655 6540
rect -4655 5620 -3655 5700
rect -3041 6540 -2041 6620
rect -3041 5700 -2961 6540
rect -2121 5700 -2041 6540
rect -3041 5620 -2041 5700
rect -1427 6540 -427 6620
rect -1427 5700 -1347 6540
rect -507 5700 -427 6540
rect -1427 5620 -427 5700
rect 187 6540 1187 6620
rect 187 5700 267 6540
rect 1107 5700 1187 6540
rect 187 5620 1187 5700
rect 1801 6540 2801 6620
rect 1801 5700 1881 6540
rect 2721 5700 2801 6540
rect 1801 5620 2801 5700
rect 3415 6540 4415 6620
rect 3415 5700 3495 6540
rect 4335 5700 4415 6540
rect 3415 5620 4415 5700
rect 5029 6540 6029 6620
rect 5029 5700 5109 6540
rect 5949 5700 6029 6540
rect 5029 5620 6029 5700
rect 6643 6540 7643 6620
rect 6643 5700 6723 6540
rect 7563 5700 7643 6540
rect 6643 5620 7643 5700
rect 8257 6540 9257 6620
rect 8257 5700 8337 6540
rect 9177 5700 9257 6540
rect 8257 5620 9257 5700
rect 9871 6540 10871 6620
rect 9871 5700 9951 6540
rect 10791 5700 10871 6540
rect 9871 5620 10871 5700
rect 11485 6540 12485 6620
rect 11485 5700 11565 6540
rect 12405 5700 12485 6540
rect 11485 5620 12485 5700
rect 13099 6540 14099 6620
rect 13099 5700 13179 6540
rect 14019 5700 14099 6540
rect 13099 5620 14099 5700
rect 14713 6540 15713 6620
rect 14713 5700 14793 6540
rect 15633 5700 15713 6540
rect 14713 5620 15713 5700
rect 16327 6540 17327 6620
rect 16327 5700 16407 6540
rect 17247 5700 17327 6540
rect 16327 5620 17327 5700
rect -17567 5180 -16567 5260
rect -17567 4340 -17487 5180
rect -16647 4340 -16567 5180
rect -17567 4260 -16567 4340
rect -15953 5180 -14953 5260
rect -15953 4340 -15873 5180
rect -15033 4340 -14953 5180
rect -15953 4260 -14953 4340
rect -14339 5180 -13339 5260
rect -14339 4340 -14259 5180
rect -13419 4340 -13339 5180
rect -14339 4260 -13339 4340
rect -12725 5180 -11725 5260
rect -12725 4340 -12645 5180
rect -11805 4340 -11725 5180
rect -12725 4260 -11725 4340
rect -11111 5180 -10111 5260
rect -11111 4340 -11031 5180
rect -10191 4340 -10111 5180
rect -11111 4260 -10111 4340
rect -9497 5180 -8497 5260
rect -9497 4340 -9417 5180
rect -8577 4340 -8497 5180
rect -9497 4260 -8497 4340
rect -7883 5180 -6883 5260
rect -7883 4340 -7803 5180
rect -6963 4340 -6883 5180
rect -7883 4260 -6883 4340
rect -6269 5180 -5269 5260
rect -6269 4340 -6189 5180
rect -5349 4340 -5269 5180
rect -6269 4260 -5269 4340
rect -4655 5180 -3655 5260
rect -4655 4340 -4575 5180
rect -3735 4340 -3655 5180
rect -4655 4260 -3655 4340
rect -3041 5180 -2041 5260
rect -3041 4340 -2961 5180
rect -2121 4340 -2041 5180
rect -3041 4260 -2041 4340
rect -1427 5180 -427 5260
rect -1427 4340 -1347 5180
rect -507 4340 -427 5180
rect -1427 4260 -427 4340
rect 187 5180 1187 5260
rect 187 4340 267 5180
rect 1107 4340 1187 5180
rect 187 4260 1187 4340
rect 1801 5180 2801 5260
rect 1801 4340 1881 5180
rect 2721 4340 2801 5180
rect 1801 4260 2801 4340
rect 3415 5180 4415 5260
rect 3415 4340 3495 5180
rect 4335 4340 4415 5180
rect 3415 4260 4415 4340
rect 5029 5180 6029 5260
rect 5029 4340 5109 5180
rect 5949 4340 6029 5180
rect 5029 4260 6029 4340
rect 6643 5180 7643 5260
rect 6643 4340 6723 5180
rect 7563 4340 7643 5180
rect 6643 4260 7643 4340
rect 8257 5180 9257 5260
rect 8257 4340 8337 5180
rect 9177 4340 9257 5180
rect 8257 4260 9257 4340
rect 9871 5180 10871 5260
rect 9871 4340 9951 5180
rect 10791 4340 10871 5180
rect 9871 4260 10871 4340
rect 11485 5180 12485 5260
rect 11485 4340 11565 5180
rect 12405 4340 12485 5180
rect 11485 4260 12485 4340
rect 13099 5180 14099 5260
rect 13099 4340 13179 5180
rect 14019 4340 14099 5180
rect 13099 4260 14099 4340
rect 14713 5180 15713 5260
rect 14713 4340 14793 5180
rect 15633 4340 15713 5180
rect 14713 4260 15713 4340
rect 16327 5180 17327 5260
rect 16327 4340 16407 5180
rect 17247 4340 17327 5180
rect 16327 4260 17327 4340
rect -17567 3820 -16567 3900
rect -17567 2980 -17487 3820
rect -16647 2980 -16567 3820
rect -17567 2900 -16567 2980
rect -15953 3820 -14953 3900
rect -15953 2980 -15873 3820
rect -15033 2980 -14953 3820
rect -15953 2900 -14953 2980
rect -14339 3820 -13339 3900
rect -14339 2980 -14259 3820
rect -13419 2980 -13339 3820
rect -14339 2900 -13339 2980
rect -12725 3820 -11725 3900
rect -12725 2980 -12645 3820
rect -11805 2980 -11725 3820
rect -12725 2900 -11725 2980
rect -11111 3820 -10111 3900
rect -11111 2980 -11031 3820
rect -10191 2980 -10111 3820
rect -11111 2900 -10111 2980
rect -9497 3820 -8497 3900
rect -9497 2980 -9417 3820
rect -8577 2980 -8497 3820
rect -9497 2900 -8497 2980
rect -7883 3820 -6883 3900
rect -7883 2980 -7803 3820
rect -6963 2980 -6883 3820
rect -7883 2900 -6883 2980
rect -6269 3820 -5269 3900
rect -6269 2980 -6189 3820
rect -5349 2980 -5269 3820
rect -6269 2900 -5269 2980
rect -4655 3820 -3655 3900
rect -4655 2980 -4575 3820
rect -3735 2980 -3655 3820
rect -4655 2900 -3655 2980
rect -3041 3820 -2041 3900
rect -3041 2980 -2961 3820
rect -2121 2980 -2041 3820
rect -3041 2900 -2041 2980
rect -1427 3820 -427 3900
rect -1427 2980 -1347 3820
rect -507 2980 -427 3820
rect -1427 2900 -427 2980
rect 187 3820 1187 3900
rect 187 2980 267 3820
rect 1107 2980 1187 3820
rect 187 2900 1187 2980
rect 1801 3820 2801 3900
rect 1801 2980 1881 3820
rect 2721 2980 2801 3820
rect 1801 2900 2801 2980
rect 3415 3820 4415 3900
rect 3415 2980 3495 3820
rect 4335 2980 4415 3820
rect 3415 2900 4415 2980
rect 5029 3820 6029 3900
rect 5029 2980 5109 3820
rect 5949 2980 6029 3820
rect 5029 2900 6029 2980
rect 6643 3820 7643 3900
rect 6643 2980 6723 3820
rect 7563 2980 7643 3820
rect 6643 2900 7643 2980
rect 8257 3820 9257 3900
rect 8257 2980 8337 3820
rect 9177 2980 9257 3820
rect 8257 2900 9257 2980
rect 9871 3820 10871 3900
rect 9871 2980 9951 3820
rect 10791 2980 10871 3820
rect 9871 2900 10871 2980
rect 11485 3820 12485 3900
rect 11485 2980 11565 3820
rect 12405 2980 12485 3820
rect 11485 2900 12485 2980
rect 13099 3820 14099 3900
rect 13099 2980 13179 3820
rect 14019 2980 14099 3820
rect 13099 2900 14099 2980
rect 14713 3820 15713 3900
rect 14713 2980 14793 3820
rect 15633 2980 15713 3820
rect 14713 2900 15713 2980
rect 16327 3820 17327 3900
rect 16327 2980 16407 3820
rect 17247 2980 17327 3820
rect 16327 2900 17327 2980
rect -17567 2460 -16567 2540
rect -17567 1620 -17487 2460
rect -16647 1620 -16567 2460
rect -17567 1540 -16567 1620
rect -15953 2460 -14953 2540
rect -15953 1620 -15873 2460
rect -15033 1620 -14953 2460
rect -15953 1540 -14953 1620
rect -14339 2460 -13339 2540
rect -14339 1620 -14259 2460
rect -13419 1620 -13339 2460
rect -14339 1540 -13339 1620
rect -12725 2460 -11725 2540
rect -12725 1620 -12645 2460
rect -11805 1620 -11725 2460
rect -12725 1540 -11725 1620
rect -11111 2460 -10111 2540
rect -11111 1620 -11031 2460
rect -10191 1620 -10111 2460
rect -11111 1540 -10111 1620
rect -9497 2460 -8497 2540
rect -9497 1620 -9417 2460
rect -8577 1620 -8497 2460
rect -9497 1540 -8497 1620
rect -7883 2460 -6883 2540
rect -7883 1620 -7803 2460
rect -6963 1620 -6883 2460
rect -7883 1540 -6883 1620
rect -6269 2460 -5269 2540
rect -6269 1620 -6189 2460
rect -5349 1620 -5269 2460
rect -6269 1540 -5269 1620
rect -4655 2460 -3655 2540
rect -4655 1620 -4575 2460
rect -3735 1620 -3655 2460
rect -4655 1540 -3655 1620
rect -3041 2460 -2041 2540
rect -3041 1620 -2961 2460
rect -2121 1620 -2041 2460
rect -3041 1540 -2041 1620
rect -1427 2460 -427 2540
rect -1427 1620 -1347 2460
rect -507 1620 -427 2460
rect -1427 1540 -427 1620
rect 187 2460 1187 2540
rect 187 1620 267 2460
rect 1107 1620 1187 2460
rect 187 1540 1187 1620
rect 1801 2460 2801 2540
rect 1801 1620 1881 2460
rect 2721 1620 2801 2460
rect 1801 1540 2801 1620
rect 3415 2460 4415 2540
rect 3415 1620 3495 2460
rect 4335 1620 4415 2460
rect 3415 1540 4415 1620
rect 5029 2460 6029 2540
rect 5029 1620 5109 2460
rect 5949 1620 6029 2460
rect 5029 1540 6029 1620
rect 6643 2460 7643 2540
rect 6643 1620 6723 2460
rect 7563 1620 7643 2460
rect 6643 1540 7643 1620
rect 8257 2460 9257 2540
rect 8257 1620 8337 2460
rect 9177 1620 9257 2460
rect 8257 1540 9257 1620
rect 9871 2460 10871 2540
rect 9871 1620 9951 2460
rect 10791 1620 10871 2460
rect 9871 1540 10871 1620
rect 11485 2460 12485 2540
rect 11485 1620 11565 2460
rect 12405 1620 12485 2460
rect 11485 1540 12485 1620
rect 13099 2460 14099 2540
rect 13099 1620 13179 2460
rect 14019 1620 14099 2460
rect 13099 1540 14099 1620
rect 14713 2460 15713 2540
rect 14713 1620 14793 2460
rect 15633 1620 15713 2460
rect 14713 1540 15713 1620
rect 16327 2460 17327 2540
rect 16327 1620 16407 2460
rect 17247 1620 17327 2460
rect 16327 1540 17327 1620
rect -17567 1100 -16567 1180
rect -17567 260 -17487 1100
rect -16647 260 -16567 1100
rect -17567 180 -16567 260
rect -15953 1100 -14953 1180
rect -15953 260 -15873 1100
rect -15033 260 -14953 1100
rect -15953 180 -14953 260
rect -14339 1100 -13339 1180
rect -14339 260 -14259 1100
rect -13419 260 -13339 1100
rect -14339 180 -13339 260
rect -12725 1100 -11725 1180
rect -12725 260 -12645 1100
rect -11805 260 -11725 1100
rect -12725 180 -11725 260
rect -11111 1100 -10111 1180
rect -11111 260 -11031 1100
rect -10191 260 -10111 1100
rect -11111 180 -10111 260
rect -9497 1100 -8497 1180
rect -9497 260 -9417 1100
rect -8577 260 -8497 1100
rect -9497 180 -8497 260
rect -7883 1100 -6883 1180
rect -7883 260 -7803 1100
rect -6963 260 -6883 1100
rect -7883 180 -6883 260
rect -6269 1100 -5269 1180
rect -6269 260 -6189 1100
rect -5349 260 -5269 1100
rect -6269 180 -5269 260
rect -4655 1100 -3655 1180
rect -4655 260 -4575 1100
rect -3735 260 -3655 1100
rect -4655 180 -3655 260
rect -3041 1100 -2041 1180
rect -3041 260 -2961 1100
rect -2121 260 -2041 1100
rect -3041 180 -2041 260
rect -1427 1100 -427 1180
rect -1427 260 -1347 1100
rect -507 260 -427 1100
rect -1427 180 -427 260
rect 187 1100 1187 1180
rect 187 260 267 1100
rect 1107 260 1187 1100
rect 187 180 1187 260
rect 1801 1100 2801 1180
rect 1801 260 1881 1100
rect 2721 260 2801 1100
rect 1801 180 2801 260
rect 3415 1100 4415 1180
rect 3415 260 3495 1100
rect 4335 260 4415 1100
rect 3415 180 4415 260
rect 5029 1100 6029 1180
rect 5029 260 5109 1100
rect 5949 260 6029 1100
rect 5029 180 6029 260
rect 6643 1100 7643 1180
rect 6643 260 6723 1100
rect 7563 260 7643 1100
rect 6643 180 7643 260
rect 8257 1100 9257 1180
rect 8257 260 8337 1100
rect 9177 260 9257 1100
rect 8257 180 9257 260
rect 9871 1100 10871 1180
rect 9871 260 9951 1100
rect 10791 260 10871 1100
rect 9871 180 10871 260
rect 11485 1100 12485 1180
rect 11485 260 11565 1100
rect 12405 260 12485 1100
rect 11485 180 12485 260
rect 13099 1100 14099 1180
rect 13099 260 13179 1100
rect 14019 260 14099 1100
rect 13099 180 14099 260
rect 14713 1100 15713 1180
rect 14713 260 14793 1100
rect 15633 260 15713 1100
rect 14713 180 15713 260
rect 16327 1100 17327 1180
rect 16327 260 16407 1100
rect 17247 260 17327 1100
rect 16327 180 17327 260
rect -17567 -260 -16567 -180
rect -17567 -1100 -17487 -260
rect -16647 -1100 -16567 -260
rect -17567 -1180 -16567 -1100
rect -15953 -260 -14953 -180
rect -15953 -1100 -15873 -260
rect -15033 -1100 -14953 -260
rect -15953 -1180 -14953 -1100
rect -14339 -260 -13339 -180
rect -14339 -1100 -14259 -260
rect -13419 -1100 -13339 -260
rect -14339 -1180 -13339 -1100
rect -12725 -260 -11725 -180
rect -12725 -1100 -12645 -260
rect -11805 -1100 -11725 -260
rect -12725 -1180 -11725 -1100
rect -11111 -260 -10111 -180
rect -11111 -1100 -11031 -260
rect -10191 -1100 -10111 -260
rect -11111 -1180 -10111 -1100
rect -9497 -260 -8497 -180
rect -9497 -1100 -9417 -260
rect -8577 -1100 -8497 -260
rect -9497 -1180 -8497 -1100
rect -7883 -260 -6883 -180
rect -7883 -1100 -7803 -260
rect -6963 -1100 -6883 -260
rect -7883 -1180 -6883 -1100
rect -6269 -260 -5269 -180
rect -6269 -1100 -6189 -260
rect -5349 -1100 -5269 -260
rect -6269 -1180 -5269 -1100
rect -4655 -260 -3655 -180
rect -4655 -1100 -4575 -260
rect -3735 -1100 -3655 -260
rect -4655 -1180 -3655 -1100
rect -3041 -260 -2041 -180
rect -3041 -1100 -2961 -260
rect -2121 -1100 -2041 -260
rect -3041 -1180 -2041 -1100
rect -1427 -260 -427 -180
rect -1427 -1100 -1347 -260
rect -507 -1100 -427 -260
rect -1427 -1180 -427 -1100
rect 187 -260 1187 -180
rect 187 -1100 267 -260
rect 1107 -1100 1187 -260
rect 187 -1180 1187 -1100
rect 1801 -260 2801 -180
rect 1801 -1100 1881 -260
rect 2721 -1100 2801 -260
rect 1801 -1180 2801 -1100
rect 3415 -260 4415 -180
rect 3415 -1100 3495 -260
rect 4335 -1100 4415 -260
rect 3415 -1180 4415 -1100
rect 5029 -260 6029 -180
rect 5029 -1100 5109 -260
rect 5949 -1100 6029 -260
rect 5029 -1180 6029 -1100
rect 6643 -260 7643 -180
rect 6643 -1100 6723 -260
rect 7563 -1100 7643 -260
rect 6643 -1180 7643 -1100
rect 8257 -260 9257 -180
rect 8257 -1100 8337 -260
rect 9177 -1100 9257 -260
rect 8257 -1180 9257 -1100
rect 9871 -260 10871 -180
rect 9871 -1100 9951 -260
rect 10791 -1100 10871 -260
rect 9871 -1180 10871 -1100
rect 11485 -260 12485 -180
rect 11485 -1100 11565 -260
rect 12405 -1100 12485 -260
rect 11485 -1180 12485 -1100
rect 13099 -260 14099 -180
rect 13099 -1100 13179 -260
rect 14019 -1100 14099 -260
rect 13099 -1180 14099 -1100
rect 14713 -260 15713 -180
rect 14713 -1100 14793 -260
rect 15633 -1100 15713 -260
rect 14713 -1180 15713 -1100
rect 16327 -260 17327 -180
rect 16327 -1100 16407 -260
rect 17247 -1100 17327 -260
rect 16327 -1180 17327 -1100
rect -17567 -1620 -16567 -1540
rect -17567 -2460 -17487 -1620
rect -16647 -2460 -16567 -1620
rect -17567 -2540 -16567 -2460
rect -15953 -1620 -14953 -1540
rect -15953 -2460 -15873 -1620
rect -15033 -2460 -14953 -1620
rect -15953 -2540 -14953 -2460
rect -14339 -1620 -13339 -1540
rect -14339 -2460 -14259 -1620
rect -13419 -2460 -13339 -1620
rect -14339 -2540 -13339 -2460
rect -12725 -1620 -11725 -1540
rect -12725 -2460 -12645 -1620
rect -11805 -2460 -11725 -1620
rect -12725 -2540 -11725 -2460
rect -11111 -1620 -10111 -1540
rect -11111 -2460 -11031 -1620
rect -10191 -2460 -10111 -1620
rect -11111 -2540 -10111 -2460
rect -9497 -1620 -8497 -1540
rect -9497 -2460 -9417 -1620
rect -8577 -2460 -8497 -1620
rect -9497 -2540 -8497 -2460
rect -7883 -1620 -6883 -1540
rect -7883 -2460 -7803 -1620
rect -6963 -2460 -6883 -1620
rect -7883 -2540 -6883 -2460
rect -6269 -1620 -5269 -1540
rect -6269 -2460 -6189 -1620
rect -5349 -2460 -5269 -1620
rect -6269 -2540 -5269 -2460
rect -4655 -1620 -3655 -1540
rect -4655 -2460 -4575 -1620
rect -3735 -2460 -3655 -1620
rect -4655 -2540 -3655 -2460
rect -3041 -1620 -2041 -1540
rect -3041 -2460 -2961 -1620
rect -2121 -2460 -2041 -1620
rect -3041 -2540 -2041 -2460
rect -1427 -1620 -427 -1540
rect -1427 -2460 -1347 -1620
rect -507 -2460 -427 -1620
rect -1427 -2540 -427 -2460
rect 187 -1620 1187 -1540
rect 187 -2460 267 -1620
rect 1107 -2460 1187 -1620
rect 187 -2540 1187 -2460
rect 1801 -1620 2801 -1540
rect 1801 -2460 1881 -1620
rect 2721 -2460 2801 -1620
rect 1801 -2540 2801 -2460
rect 3415 -1620 4415 -1540
rect 3415 -2460 3495 -1620
rect 4335 -2460 4415 -1620
rect 3415 -2540 4415 -2460
rect 5029 -1620 6029 -1540
rect 5029 -2460 5109 -1620
rect 5949 -2460 6029 -1620
rect 5029 -2540 6029 -2460
rect 6643 -1620 7643 -1540
rect 6643 -2460 6723 -1620
rect 7563 -2460 7643 -1620
rect 6643 -2540 7643 -2460
rect 8257 -1620 9257 -1540
rect 8257 -2460 8337 -1620
rect 9177 -2460 9257 -1620
rect 8257 -2540 9257 -2460
rect 9871 -1620 10871 -1540
rect 9871 -2460 9951 -1620
rect 10791 -2460 10871 -1620
rect 9871 -2540 10871 -2460
rect 11485 -1620 12485 -1540
rect 11485 -2460 11565 -1620
rect 12405 -2460 12485 -1620
rect 11485 -2540 12485 -2460
rect 13099 -1620 14099 -1540
rect 13099 -2460 13179 -1620
rect 14019 -2460 14099 -1620
rect 13099 -2540 14099 -2460
rect 14713 -1620 15713 -1540
rect 14713 -2460 14793 -1620
rect 15633 -2460 15713 -1620
rect 14713 -2540 15713 -2460
rect 16327 -1620 17327 -1540
rect 16327 -2460 16407 -1620
rect 17247 -2460 17327 -1620
rect 16327 -2540 17327 -2460
rect -17567 -2980 -16567 -2900
rect -17567 -3820 -17487 -2980
rect -16647 -3820 -16567 -2980
rect -17567 -3900 -16567 -3820
rect -15953 -2980 -14953 -2900
rect -15953 -3820 -15873 -2980
rect -15033 -3820 -14953 -2980
rect -15953 -3900 -14953 -3820
rect -14339 -2980 -13339 -2900
rect -14339 -3820 -14259 -2980
rect -13419 -3820 -13339 -2980
rect -14339 -3900 -13339 -3820
rect -12725 -2980 -11725 -2900
rect -12725 -3820 -12645 -2980
rect -11805 -3820 -11725 -2980
rect -12725 -3900 -11725 -3820
rect -11111 -2980 -10111 -2900
rect -11111 -3820 -11031 -2980
rect -10191 -3820 -10111 -2980
rect -11111 -3900 -10111 -3820
rect -9497 -2980 -8497 -2900
rect -9497 -3820 -9417 -2980
rect -8577 -3820 -8497 -2980
rect -9497 -3900 -8497 -3820
rect -7883 -2980 -6883 -2900
rect -7883 -3820 -7803 -2980
rect -6963 -3820 -6883 -2980
rect -7883 -3900 -6883 -3820
rect -6269 -2980 -5269 -2900
rect -6269 -3820 -6189 -2980
rect -5349 -3820 -5269 -2980
rect -6269 -3900 -5269 -3820
rect -4655 -2980 -3655 -2900
rect -4655 -3820 -4575 -2980
rect -3735 -3820 -3655 -2980
rect -4655 -3900 -3655 -3820
rect -3041 -2980 -2041 -2900
rect -3041 -3820 -2961 -2980
rect -2121 -3820 -2041 -2980
rect -3041 -3900 -2041 -3820
rect -1427 -2980 -427 -2900
rect -1427 -3820 -1347 -2980
rect -507 -3820 -427 -2980
rect -1427 -3900 -427 -3820
rect 187 -2980 1187 -2900
rect 187 -3820 267 -2980
rect 1107 -3820 1187 -2980
rect 187 -3900 1187 -3820
rect 1801 -2980 2801 -2900
rect 1801 -3820 1881 -2980
rect 2721 -3820 2801 -2980
rect 1801 -3900 2801 -3820
rect 3415 -2980 4415 -2900
rect 3415 -3820 3495 -2980
rect 4335 -3820 4415 -2980
rect 3415 -3900 4415 -3820
rect 5029 -2980 6029 -2900
rect 5029 -3820 5109 -2980
rect 5949 -3820 6029 -2980
rect 5029 -3900 6029 -3820
rect 6643 -2980 7643 -2900
rect 6643 -3820 6723 -2980
rect 7563 -3820 7643 -2980
rect 6643 -3900 7643 -3820
rect 8257 -2980 9257 -2900
rect 8257 -3820 8337 -2980
rect 9177 -3820 9257 -2980
rect 8257 -3900 9257 -3820
rect 9871 -2980 10871 -2900
rect 9871 -3820 9951 -2980
rect 10791 -3820 10871 -2980
rect 9871 -3900 10871 -3820
rect 11485 -2980 12485 -2900
rect 11485 -3820 11565 -2980
rect 12405 -3820 12485 -2980
rect 11485 -3900 12485 -3820
rect 13099 -2980 14099 -2900
rect 13099 -3820 13179 -2980
rect 14019 -3820 14099 -2980
rect 13099 -3900 14099 -3820
rect 14713 -2980 15713 -2900
rect 14713 -3820 14793 -2980
rect 15633 -3820 15713 -2980
rect 14713 -3900 15713 -3820
rect 16327 -2980 17327 -2900
rect 16327 -3820 16407 -2980
rect 17247 -3820 17327 -2980
rect 16327 -3900 17327 -3820
rect -17567 -4340 -16567 -4260
rect -17567 -5180 -17487 -4340
rect -16647 -5180 -16567 -4340
rect -17567 -5260 -16567 -5180
rect -15953 -4340 -14953 -4260
rect -15953 -5180 -15873 -4340
rect -15033 -5180 -14953 -4340
rect -15953 -5260 -14953 -5180
rect -14339 -4340 -13339 -4260
rect -14339 -5180 -14259 -4340
rect -13419 -5180 -13339 -4340
rect -14339 -5260 -13339 -5180
rect -12725 -4340 -11725 -4260
rect -12725 -5180 -12645 -4340
rect -11805 -5180 -11725 -4340
rect -12725 -5260 -11725 -5180
rect -11111 -4340 -10111 -4260
rect -11111 -5180 -11031 -4340
rect -10191 -5180 -10111 -4340
rect -11111 -5260 -10111 -5180
rect -9497 -4340 -8497 -4260
rect -9497 -5180 -9417 -4340
rect -8577 -5180 -8497 -4340
rect -9497 -5260 -8497 -5180
rect -7883 -4340 -6883 -4260
rect -7883 -5180 -7803 -4340
rect -6963 -5180 -6883 -4340
rect -7883 -5260 -6883 -5180
rect -6269 -4340 -5269 -4260
rect -6269 -5180 -6189 -4340
rect -5349 -5180 -5269 -4340
rect -6269 -5260 -5269 -5180
rect -4655 -4340 -3655 -4260
rect -4655 -5180 -4575 -4340
rect -3735 -5180 -3655 -4340
rect -4655 -5260 -3655 -5180
rect -3041 -4340 -2041 -4260
rect -3041 -5180 -2961 -4340
rect -2121 -5180 -2041 -4340
rect -3041 -5260 -2041 -5180
rect -1427 -4340 -427 -4260
rect -1427 -5180 -1347 -4340
rect -507 -5180 -427 -4340
rect -1427 -5260 -427 -5180
rect 187 -4340 1187 -4260
rect 187 -5180 267 -4340
rect 1107 -5180 1187 -4340
rect 187 -5260 1187 -5180
rect 1801 -4340 2801 -4260
rect 1801 -5180 1881 -4340
rect 2721 -5180 2801 -4340
rect 1801 -5260 2801 -5180
rect 3415 -4340 4415 -4260
rect 3415 -5180 3495 -4340
rect 4335 -5180 4415 -4340
rect 3415 -5260 4415 -5180
rect 5029 -4340 6029 -4260
rect 5029 -5180 5109 -4340
rect 5949 -5180 6029 -4340
rect 5029 -5260 6029 -5180
rect 6643 -4340 7643 -4260
rect 6643 -5180 6723 -4340
rect 7563 -5180 7643 -4340
rect 6643 -5260 7643 -5180
rect 8257 -4340 9257 -4260
rect 8257 -5180 8337 -4340
rect 9177 -5180 9257 -4340
rect 8257 -5260 9257 -5180
rect 9871 -4340 10871 -4260
rect 9871 -5180 9951 -4340
rect 10791 -5180 10871 -4340
rect 9871 -5260 10871 -5180
rect 11485 -4340 12485 -4260
rect 11485 -5180 11565 -4340
rect 12405 -5180 12485 -4340
rect 11485 -5260 12485 -5180
rect 13099 -4340 14099 -4260
rect 13099 -5180 13179 -4340
rect 14019 -5180 14099 -4340
rect 13099 -5260 14099 -5180
rect 14713 -4340 15713 -4260
rect 14713 -5180 14793 -4340
rect 15633 -5180 15713 -4340
rect 14713 -5260 15713 -5180
rect 16327 -4340 17327 -4260
rect 16327 -5180 16407 -4340
rect 17247 -5180 17327 -4340
rect 16327 -5260 17327 -5180
rect -17567 -5700 -16567 -5620
rect -17567 -6540 -17487 -5700
rect -16647 -6540 -16567 -5700
rect -17567 -6620 -16567 -6540
rect -15953 -5700 -14953 -5620
rect -15953 -6540 -15873 -5700
rect -15033 -6540 -14953 -5700
rect -15953 -6620 -14953 -6540
rect -14339 -5700 -13339 -5620
rect -14339 -6540 -14259 -5700
rect -13419 -6540 -13339 -5700
rect -14339 -6620 -13339 -6540
rect -12725 -5700 -11725 -5620
rect -12725 -6540 -12645 -5700
rect -11805 -6540 -11725 -5700
rect -12725 -6620 -11725 -6540
rect -11111 -5700 -10111 -5620
rect -11111 -6540 -11031 -5700
rect -10191 -6540 -10111 -5700
rect -11111 -6620 -10111 -6540
rect -9497 -5700 -8497 -5620
rect -9497 -6540 -9417 -5700
rect -8577 -6540 -8497 -5700
rect -9497 -6620 -8497 -6540
rect -7883 -5700 -6883 -5620
rect -7883 -6540 -7803 -5700
rect -6963 -6540 -6883 -5700
rect -7883 -6620 -6883 -6540
rect -6269 -5700 -5269 -5620
rect -6269 -6540 -6189 -5700
rect -5349 -6540 -5269 -5700
rect -6269 -6620 -5269 -6540
rect -4655 -5700 -3655 -5620
rect -4655 -6540 -4575 -5700
rect -3735 -6540 -3655 -5700
rect -4655 -6620 -3655 -6540
rect -3041 -5700 -2041 -5620
rect -3041 -6540 -2961 -5700
rect -2121 -6540 -2041 -5700
rect -3041 -6620 -2041 -6540
rect -1427 -5700 -427 -5620
rect -1427 -6540 -1347 -5700
rect -507 -6540 -427 -5700
rect -1427 -6620 -427 -6540
rect 187 -5700 1187 -5620
rect 187 -6540 267 -5700
rect 1107 -6540 1187 -5700
rect 187 -6620 1187 -6540
rect 1801 -5700 2801 -5620
rect 1801 -6540 1881 -5700
rect 2721 -6540 2801 -5700
rect 1801 -6620 2801 -6540
rect 3415 -5700 4415 -5620
rect 3415 -6540 3495 -5700
rect 4335 -6540 4415 -5700
rect 3415 -6620 4415 -6540
rect 5029 -5700 6029 -5620
rect 5029 -6540 5109 -5700
rect 5949 -6540 6029 -5700
rect 5029 -6620 6029 -6540
rect 6643 -5700 7643 -5620
rect 6643 -6540 6723 -5700
rect 7563 -6540 7643 -5700
rect 6643 -6620 7643 -6540
rect 8257 -5700 9257 -5620
rect 8257 -6540 8337 -5700
rect 9177 -6540 9257 -5700
rect 8257 -6620 9257 -6540
rect 9871 -5700 10871 -5620
rect 9871 -6540 9951 -5700
rect 10791 -6540 10871 -5700
rect 9871 -6620 10871 -6540
rect 11485 -5700 12485 -5620
rect 11485 -6540 11565 -5700
rect 12405 -6540 12485 -5700
rect 11485 -6620 12485 -6540
rect 13099 -5700 14099 -5620
rect 13099 -6540 13179 -5700
rect 14019 -6540 14099 -5700
rect 13099 -6620 14099 -6540
rect 14713 -5700 15713 -5620
rect 14713 -6540 14793 -5700
rect 15633 -6540 15713 -5700
rect 14713 -6620 15713 -6540
rect 16327 -5700 17327 -5620
rect 16327 -6540 16407 -5700
rect 17247 -6540 17327 -5700
rect 16327 -6620 17327 -6540
rect -17567 -7060 -16567 -6980
rect -17567 -7900 -17487 -7060
rect -16647 -7900 -16567 -7060
rect -17567 -7980 -16567 -7900
rect -15953 -7060 -14953 -6980
rect -15953 -7900 -15873 -7060
rect -15033 -7900 -14953 -7060
rect -15953 -7980 -14953 -7900
rect -14339 -7060 -13339 -6980
rect -14339 -7900 -14259 -7060
rect -13419 -7900 -13339 -7060
rect -14339 -7980 -13339 -7900
rect -12725 -7060 -11725 -6980
rect -12725 -7900 -12645 -7060
rect -11805 -7900 -11725 -7060
rect -12725 -7980 -11725 -7900
rect -11111 -7060 -10111 -6980
rect -11111 -7900 -11031 -7060
rect -10191 -7900 -10111 -7060
rect -11111 -7980 -10111 -7900
rect -9497 -7060 -8497 -6980
rect -9497 -7900 -9417 -7060
rect -8577 -7900 -8497 -7060
rect -9497 -7980 -8497 -7900
rect -7883 -7060 -6883 -6980
rect -7883 -7900 -7803 -7060
rect -6963 -7900 -6883 -7060
rect -7883 -7980 -6883 -7900
rect -6269 -7060 -5269 -6980
rect -6269 -7900 -6189 -7060
rect -5349 -7900 -5269 -7060
rect -6269 -7980 -5269 -7900
rect -4655 -7060 -3655 -6980
rect -4655 -7900 -4575 -7060
rect -3735 -7900 -3655 -7060
rect -4655 -7980 -3655 -7900
rect -3041 -7060 -2041 -6980
rect -3041 -7900 -2961 -7060
rect -2121 -7900 -2041 -7060
rect -3041 -7980 -2041 -7900
rect -1427 -7060 -427 -6980
rect -1427 -7900 -1347 -7060
rect -507 -7900 -427 -7060
rect -1427 -7980 -427 -7900
rect 187 -7060 1187 -6980
rect 187 -7900 267 -7060
rect 1107 -7900 1187 -7060
rect 187 -7980 1187 -7900
rect 1801 -7060 2801 -6980
rect 1801 -7900 1881 -7060
rect 2721 -7900 2801 -7060
rect 1801 -7980 2801 -7900
rect 3415 -7060 4415 -6980
rect 3415 -7900 3495 -7060
rect 4335 -7900 4415 -7060
rect 3415 -7980 4415 -7900
rect 5029 -7060 6029 -6980
rect 5029 -7900 5109 -7060
rect 5949 -7900 6029 -7060
rect 5029 -7980 6029 -7900
rect 6643 -7060 7643 -6980
rect 6643 -7900 6723 -7060
rect 7563 -7900 7643 -7060
rect 6643 -7980 7643 -7900
rect 8257 -7060 9257 -6980
rect 8257 -7900 8337 -7060
rect 9177 -7900 9257 -7060
rect 8257 -7980 9257 -7900
rect 9871 -7060 10871 -6980
rect 9871 -7900 9951 -7060
rect 10791 -7900 10871 -7060
rect 9871 -7980 10871 -7900
rect 11485 -7060 12485 -6980
rect 11485 -7900 11565 -7060
rect 12405 -7900 12485 -7060
rect 11485 -7980 12485 -7900
rect 13099 -7060 14099 -6980
rect 13099 -7900 13179 -7060
rect 14019 -7900 14099 -7060
rect 13099 -7980 14099 -7900
rect 14713 -7060 15713 -6980
rect 14713 -7900 14793 -7060
rect 15633 -7900 15713 -7060
rect 14713 -7980 15713 -7900
rect 16327 -7060 17327 -6980
rect 16327 -7900 16407 -7060
rect 17247 -7900 17327 -7060
rect 16327 -7980 17327 -7900
<< mimcapcontact >>
rect -17487 7060 -16647 7900
rect -15873 7060 -15033 7900
rect -14259 7060 -13419 7900
rect -12645 7060 -11805 7900
rect -11031 7060 -10191 7900
rect -9417 7060 -8577 7900
rect -7803 7060 -6963 7900
rect -6189 7060 -5349 7900
rect -4575 7060 -3735 7900
rect -2961 7060 -2121 7900
rect -1347 7060 -507 7900
rect 267 7060 1107 7900
rect 1881 7060 2721 7900
rect 3495 7060 4335 7900
rect 5109 7060 5949 7900
rect 6723 7060 7563 7900
rect 8337 7060 9177 7900
rect 9951 7060 10791 7900
rect 11565 7060 12405 7900
rect 13179 7060 14019 7900
rect 14793 7060 15633 7900
rect 16407 7060 17247 7900
rect -17487 5700 -16647 6540
rect -15873 5700 -15033 6540
rect -14259 5700 -13419 6540
rect -12645 5700 -11805 6540
rect -11031 5700 -10191 6540
rect -9417 5700 -8577 6540
rect -7803 5700 -6963 6540
rect -6189 5700 -5349 6540
rect -4575 5700 -3735 6540
rect -2961 5700 -2121 6540
rect -1347 5700 -507 6540
rect 267 5700 1107 6540
rect 1881 5700 2721 6540
rect 3495 5700 4335 6540
rect 5109 5700 5949 6540
rect 6723 5700 7563 6540
rect 8337 5700 9177 6540
rect 9951 5700 10791 6540
rect 11565 5700 12405 6540
rect 13179 5700 14019 6540
rect 14793 5700 15633 6540
rect 16407 5700 17247 6540
rect -17487 4340 -16647 5180
rect -15873 4340 -15033 5180
rect -14259 4340 -13419 5180
rect -12645 4340 -11805 5180
rect -11031 4340 -10191 5180
rect -9417 4340 -8577 5180
rect -7803 4340 -6963 5180
rect -6189 4340 -5349 5180
rect -4575 4340 -3735 5180
rect -2961 4340 -2121 5180
rect -1347 4340 -507 5180
rect 267 4340 1107 5180
rect 1881 4340 2721 5180
rect 3495 4340 4335 5180
rect 5109 4340 5949 5180
rect 6723 4340 7563 5180
rect 8337 4340 9177 5180
rect 9951 4340 10791 5180
rect 11565 4340 12405 5180
rect 13179 4340 14019 5180
rect 14793 4340 15633 5180
rect 16407 4340 17247 5180
rect -17487 2980 -16647 3820
rect -15873 2980 -15033 3820
rect -14259 2980 -13419 3820
rect -12645 2980 -11805 3820
rect -11031 2980 -10191 3820
rect -9417 2980 -8577 3820
rect -7803 2980 -6963 3820
rect -6189 2980 -5349 3820
rect -4575 2980 -3735 3820
rect -2961 2980 -2121 3820
rect -1347 2980 -507 3820
rect 267 2980 1107 3820
rect 1881 2980 2721 3820
rect 3495 2980 4335 3820
rect 5109 2980 5949 3820
rect 6723 2980 7563 3820
rect 8337 2980 9177 3820
rect 9951 2980 10791 3820
rect 11565 2980 12405 3820
rect 13179 2980 14019 3820
rect 14793 2980 15633 3820
rect 16407 2980 17247 3820
rect -17487 1620 -16647 2460
rect -15873 1620 -15033 2460
rect -14259 1620 -13419 2460
rect -12645 1620 -11805 2460
rect -11031 1620 -10191 2460
rect -9417 1620 -8577 2460
rect -7803 1620 -6963 2460
rect -6189 1620 -5349 2460
rect -4575 1620 -3735 2460
rect -2961 1620 -2121 2460
rect -1347 1620 -507 2460
rect 267 1620 1107 2460
rect 1881 1620 2721 2460
rect 3495 1620 4335 2460
rect 5109 1620 5949 2460
rect 6723 1620 7563 2460
rect 8337 1620 9177 2460
rect 9951 1620 10791 2460
rect 11565 1620 12405 2460
rect 13179 1620 14019 2460
rect 14793 1620 15633 2460
rect 16407 1620 17247 2460
rect -17487 260 -16647 1100
rect -15873 260 -15033 1100
rect -14259 260 -13419 1100
rect -12645 260 -11805 1100
rect -11031 260 -10191 1100
rect -9417 260 -8577 1100
rect -7803 260 -6963 1100
rect -6189 260 -5349 1100
rect -4575 260 -3735 1100
rect -2961 260 -2121 1100
rect -1347 260 -507 1100
rect 267 260 1107 1100
rect 1881 260 2721 1100
rect 3495 260 4335 1100
rect 5109 260 5949 1100
rect 6723 260 7563 1100
rect 8337 260 9177 1100
rect 9951 260 10791 1100
rect 11565 260 12405 1100
rect 13179 260 14019 1100
rect 14793 260 15633 1100
rect 16407 260 17247 1100
rect -17487 -1100 -16647 -260
rect -15873 -1100 -15033 -260
rect -14259 -1100 -13419 -260
rect -12645 -1100 -11805 -260
rect -11031 -1100 -10191 -260
rect -9417 -1100 -8577 -260
rect -7803 -1100 -6963 -260
rect -6189 -1100 -5349 -260
rect -4575 -1100 -3735 -260
rect -2961 -1100 -2121 -260
rect -1347 -1100 -507 -260
rect 267 -1100 1107 -260
rect 1881 -1100 2721 -260
rect 3495 -1100 4335 -260
rect 5109 -1100 5949 -260
rect 6723 -1100 7563 -260
rect 8337 -1100 9177 -260
rect 9951 -1100 10791 -260
rect 11565 -1100 12405 -260
rect 13179 -1100 14019 -260
rect 14793 -1100 15633 -260
rect 16407 -1100 17247 -260
rect -17487 -2460 -16647 -1620
rect -15873 -2460 -15033 -1620
rect -14259 -2460 -13419 -1620
rect -12645 -2460 -11805 -1620
rect -11031 -2460 -10191 -1620
rect -9417 -2460 -8577 -1620
rect -7803 -2460 -6963 -1620
rect -6189 -2460 -5349 -1620
rect -4575 -2460 -3735 -1620
rect -2961 -2460 -2121 -1620
rect -1347 -2460 -507 -1620
rect 267 -2460 1107 -1620
rect 1881 -2460 2721 -1620
rect 3495 -2460 4335 -1620
rect 5109 -2460 5949 -1620
rect 6723 -2460 7563 -1620
rect 8337 -2460 9177 -1620
rect 9951 -2460 10791 -1620
rect 11565 -2460 12405 -1620
rect 13179 -2460 14019 -1620
rect 14793 -2460 15633 -1620
rect 16407 -2460 17247 -1620
rect -17487 -3820 -16647 -2980
rect -15873 -3820 -15033 -2980
rect -14259 -3820 -13419 -2980
rect -12645 -3820 -11805 -2980
rect -11031 -3820 -10191 -2980
rect -9417 -3820 -8577 -2980
rect -7803 -3820 -6963 -2980
rect -6189 -3820 -5349 -2980
rect -4575 -3820 -3735 -2980
rect -2961 -3820 -2121 -2980
rect -1347 -3820 -507 -2980
rect 267 -3820 1107 -2980
rect 1881 -3820 2721 -2980
rect 3495 -3820 4335 -2980
rect 5109 -3820 5949 -2980
rect 6723 -3820 7563 -2980
rect 8337 -3820 9177 -2980
rect 9951 -3820 10791 -2980
rect 11565 -3820 12405 -2980
rect 13179 -3820 14019 -2980
rect 14793 -3820 15633 -2980
rect 16407 -3820 17247 -2980
rect -17487 -5180 -16647 -4340
rect -15873 -5180 -15033 -4340
rect -14259 -5180 -13419 -4340
rect -12645 -5180 -11805 -4340
rect -11031 -5180 -10191 -4340
rect -9417 -5180 -8577 -4340
rect -7803 -5180 -6963 -4340
rect -6189 -5180 -5349 -4340
rect -4575 -5180 -3735 -4340
rect -2961 -5180 -2121 -4340
rect -1347 -5180 -507 -4340
rect 267 -5180 1107 -4340
rect 1881 -5180 2721 -4340
rect 3495 -5180 4335 -4340
rect 5109 -5180 5949 -4340
rect 6723 -5180 7563 -4340
rect 8337 -5180 9177 -4340
rect 9951 -5180 10791 -4340
rect 11565 -5180 12405 -4340
rect 13179 -5180 14019 -4340
rect 14793 -5180 15633 -4340
rect 16407 -5180 17247 -4340
rect -17487 -6540 -16647 -5700
rect -15873 -6540 -15033 -5700
rect -14259 -6540 -13419 -5700
rect -12645 -6540 -11805 -5700
rect -11031 -6540 -10191 -5700
rect -9417 -6540 -8577 -5700
rect -7803 -6540 -6963 -5700
rect -6189 -6540 -5349 -5700
rect -4575 -6540 -3735 -5700
rect -2961 -6540 -2121 -5700
rect -1347 -6540 -507 -5700
rect 267 -6540 1107 -5700
rect 1881 -6540 2721 -5700
rect 3495 -6540 4335 -5700
rect 5109 -6540 5949 -5700
rect 6723 -6540 7563 -5700
rect 8337 -6540 9177 -5700
rect 9951 -6540 10791 -5700
rect 11565 -6540 12405 -5700
rect 13179 -6540 14019 -5700
rect 14793 -6540 15633 -5700
rect 16407 -6540 17247 -5700
rect -17487 -7900 -16647 -7060
rect -15873 -7900 -15033 -7060
rect -14259 -7900 -13419 -7060
rect -12645 -7900 -11805 -7060
rect -11031 -7900 -10191 -7060
rect -9417 -7900 -8577 -7060
rect -7803 -7900 -6963 -7060
rect -6189 -7900 -5349 -7060
rect -4575 -7900 -3735 -7060
rect -2961 -7900 -2121 -7060
rect -1347 -7900 -507 -7060
rect 267 -7900 1107 -7060
rect 1881 -7900 2721 -7060
rect 3495 -7900 4335 -7060
rect 5109 -7900 5949 -7060
rect 6723 -7900 7563 -7060
rect 8337 -7900 9177 -7060
rect 9951 -7900 10791 -7060
rect 11565 -7900 12405 -7060
rect 13179 -7900 14019 -7060
rect 14793 -7900 15633 -7060
rect 16407 -7900 17247 -7060
<< metal4 >>
rect -17687 8033 -16207 8100
rect -17687 7980 -16357 8033
rect -17687 6980 -17567 7980
rect -16567 6980 -16357 7980
rect -17687 6927 -16357 6980
rect -16269 6927 -16207 8033
rect -17687 6860 -16207 6927
rect -16073 8033 -14593 8100
rect -16073 7980 -14743 8033
rect -16073 6980 -15953 7980
rect -14953 6980 -14743 7980
rect -16073 6927 -14743 6980
rect -14655 6927 -14593 8033
rect -16073 6860 -14593 6927
rect -14459 8033 -12979 8100
rect -14459 7980 -13129 8033
rect -14459 6980 -14339 7980
rect -13339 6980 -13129 7980
rect -14459 6927 -13129 6980
rect -13041 6927 -12979 8033
rect -14459 6860 -12979 6927
rect -12845 8033 -11365 8100
rect -12845 7980 -11515 8033
rect -12845 6980 -12725 7980
rect -11725 6980 -11515 7980
rect -12845 6927 -11515 6980
rect -11427 6927 -11365 8033
rect -12845 6860 -11365 6927
rect -11231 8033 -9751 8100
rect -11231 7980 -9901 8033
rect -11231 6980 -11111 7980
rect -10111 6980 -9901 7980
rect -11231 6927 -9901 6980
rect -9813 6927 -9751 8033
rect -11231 6860 -9751 6927
rect -9617 8033 -8137 8100
rect -9617 7980 -8287 8033
rect -9617 6980 -9497 7980
rect -8497 6980 -8287 7980
rect -9617 6927 -8287 6980
rect -8199 6927 -8137 8033
rect -9617 6860 -8137 6927
rect -8003 8033 -6523 8100
rect -8003 7980 -6673 8033
rect -8003 6980 -7883 7980
rect -6883 6980 -6673 7980
rect -8003 6927 -6673 6980
rect -6585 6927 -6523 8033
rect -8003 6860 -6523 6927
rect -6389 8033 -4909 8100
rect -6389 7980 -5059 8033
rect -6389 6980 -6269 7980
rect -5269 6980 -5059 7980
rect -6389 6927 -5059 6980
rect -4971 6927 -4909 8033
rect -6389 6860 -4909 6927
rect -4775 8033 -3295 8100
rect -4775 7980 -3445 8033
rect -4775 6980 -4655 7980
rect -3655 6980 -3445 7980
rect -4775 6927 -3445 6980
rect -3357 6927 -3295 8033
rect -4775 6860 -3295 6927
rect -3161 8033 -1681 8100
rect -3161 7980 -1831 8033
rect -3161 6980 -3041 7980
rect -2041 6980 -1831 7980
rect -3161 6927 -1831 6980
rect -1743 6927 -1681 8033
rect -3161 6860 -1681 6927
rect -1547 8033 -67 8100
rect -1547 7980 -217 8033
rect -1547 6980 -1427 7980
rect -427 6980 -217 7980
rect -1547 6927 -217 6980
rect -129 6927 -67 8033
rect -1547 6860 -67 6927
rect 67 8033 1547 8100
rect 67 7980 1397 8033
rect 67 6980 187 7980
rect 1187 6980 1397 7980
rect 67 6927 1397 6980
rect 1485 6927 1547 8033
rect 67 6860 1547 6927
rect 1681 8033 3161 8100
rect 1681 7980 3011 8033
rect 1681 6980 1801 7980
rect 2801 6980 3011 7980
rect 1681 6927 3011 6980
rect 3099 6927 3161 8033
rect 1681 6860 3161 6927
rect 3295 8033 4775 8100
rect 3295 7980 4625 8033
rect 3295 6980 3415 7980
rect 4415 6980 4625 7980
rect 3295 6927 4625 6980
rect 4713 6927 4775 8033
rect 3295 6860 4775 6927
rect 4909 8033 6389 8100
rect 4909 7980 6239 8033
rect 4909 6980 5029 7980
rect 6029 6980 6239 7980
rect 4909 6927 6239 6980
rect 6327 6927 6389 8033
rect 4909 6860 6389 6927
rect 6523 8033 8003 8100
rect 6523 7980 7853 8033
rect 6523 6980 6643 7980
rect 7643 6980 7853 7980
rect 6523 6927 7853 6980
rect 7941 6927 8003 8033
rect 6523 6860 8003 6927
rect 8137 8033 9617 8100
rect 8137 7980 9467 8033
rect 8137 6980 8257 7980
rect 9257 6980 9467 7980
rect 8137 6927 9467 6980
rect 9555 6927 9617 8033
rect 8137 6860 9617 6927
rect 9751 8033 11231 8100
rect 9751 7980 11081 8033
rect 9751 6980 9871 7980
rect 10871 6980 11081 7980
rect 9751 6927 11081 6980
rect 11169 6927 11231 8033
rect 9751 6860 11231 6927
rect 11365 8033 12845 8100
rect 11365 7980 12695 8033
rect 11365 6980 11485 7980
rect 12485 6980 12695 7980
rect 11365 6927 12695 6980
rect 12783 6927 12845 8033
rect 11365 6860 12845 6927
rect 12979 8033 14459 8100
rect 12979 7980 14309 8033
rect 12979 6980 13099 7980
rect 14099 6980 14309 7980
rect 12979 6927 14309 6980
rect 14397 6927 14459 8033
rect 12979 6860 14459 6927
rect 14593 8033 16073 8100
rect 14593 7980 15923 8033
rect 14593 6980 14713 7980
rect 15713 6980 15923 7980
rect 14593 6927 15923 6980
rect 16011 6927 16073 8033
rect 14593 6860 16073 6927
rect 16207 8033 17687 8100
rect 16207 7980 17537 8033
rect 16207 6980 16327 7980
rect 17327 6980 17537 7980
rect 16207 6927 17537 6980
rect 17625 6927 17687 8033
rect 16207 6860 17687 6927
rect -17687 6673 -16207 6740
rect -17687 6620 -16357 6673
rect -17687 5620 -17567 6620
rect -16567 5620 -16357 6620
rect -17687 5567 -16357 5620
rect -16269 5567 -16207 6673
rect -17687 5500 -16207 5567
rect -16073 6673 -14593 6740
rect -16073 6620 -14743 6673
rect -16073 5620 -15953 6620
rect -14953 5620 -14743 6620
rect -16073 5567 -14743 5620
rect -14655 5567 -14593 6673
rect -16073 5500 -14593 5567
rect -14459 6673 -12979 6740
rect -14459 6620 -13129 6673
rect -14459 5620 -14339 6620
rect -13339 5620 -13129 6620
rect -14459 5567 -13129 5620
rect -13041 5567 -12979 6673
rect -14459 5500 -12979 5567
rect -12845 6673 -11365 6740
rect -12845 6620 -11515 6673
rect -12845 5620 -12725 6620
rect -11725 5620 -11515 6620
rect -12845 5567 -11515 5620
rect -11427 5567 -11365 6673
rect -12845 5500 -11365 5567
rect -11231 6673 -9751 6740
rect -11231 6620 -9901 6673
rect -11231 5620 -11111 6620
rect -10111 5620 -9901 6620
rect -11231 5567 -9901 5620
rect -9813 5567 -9751 6673
rect -11231 5500 -9751 5567
rect -9617 6673 -8137 6740
rect -9617 6620 -8287 6673
rect -9617 5620 -9497 6620
rect -8497 5620 -8287 6620
rect -9617 5567 -8287 5620
rect -8199 5567 -8137 6673
rect -9617 5500 -8137 5567
rect -8003 6673 -6523 6740
rect -8003 6620 -6673 6673
rect -8003 5620 -7883 6620
rect -6883 5620 -6673 6620
rect -8003 5567 -6673 5620
rect -6585 5567 -6523 6673
rect -8003 5500 -6523 5567
rect -6389 6673 -4909 6740
rect -6389 6620 -5059 6673
rect -6389 5620 -6269 6620
rect -5269 5620 -5059 6620
rect -6389 5567 -5059 5620
rect -4971 5567 -4909 6673
rect -6389 5500 -4909 5567
rect -4775 6673 -3295 6740
rect -4775 6620 -3445 6673
rect -4775 5620 -4655 6620
rect -3655 5620 -3445 6620
rect -4775 5567 -3445 5620
rect -3357 5567 -3295 6673
rect -4775 5500 -3295 5567
rect -3161 6673 -1681 6740
rect -3161 6620 -1831 6673
rect -3161 5620 -3041 6620
rect -2041 5620 -1831 6620
rect -3161 5567 -1831 5620
rect -1743 5567 -1681 6673
rect -3161 5500 -1681 5567
rect -1547 6673 -67 6740
rect -1547 6620 -217 6673
rect -1547 5620 -1427 6620
rect -427 5620 -217 6620
rect -1547 5567 -217 5620
rect -129 5567 -67 6673
rect -1547 5500 -67 5567
rect 67 6673 1547 6740
rect 67 6620 1397 6673
rect 67 5620 187 6620
rect 1187 5620 1397 6620
rect 67 5567 1397 5620
rect 1485 5567 1547 6673
rect 67 5500 1547 5567
rect 1681 6673 3161 6740
rect 1681 6620 3011 6673
rect 1681 5620 1801 6620
rect 2801 5620 3011 6620
rect 1681 5567 3011 5620
rect 3099 5567 3161 6673
rect 1681 5500 3161 5567
rect 3295 6673 4775 6740
rect 3295 6620 4625 6673
rect 3295 5620 3415 6620
rect 4415 5620 4625 6620
rect 3295 5567 4625 5620
rect 4713 5567 4775 6673
rect 3295 5500 4775 5567
rect 4909 6673 6389 6740
rect 4909 6620 6239 6673
rect 4909 5620 5029 6620
rect 6029 5620 6239 6620
rect 4909 5567 6239 5620
rect 6327 5567 6389 6673
rect 4909 5500 6389 5567
rect 6523 6673 8003 6740
rect 6523 6620 7853 6673
rect 6523 5620 6643 6620
rect 7643 5620 7853 6620
rect 6523 5567 7853 5620
rect 7941 5567 8003 6673
rect 6523 5500 8003 5567
rect 8137 6673 9617 6740
rect 8137 6620 9467 6673
rect 8137 5620 8257 6620
rect 9257 5620 9467 6620
rect 8137 5567 9467 5620
rect 9555 5567 9617 6673
rect 8137 5500 9617 5567
rect 9751 6673 11231 6740
rect 9751 6620 11081 6673
rect 9751 5620 9871 6620
rect 10871 5620 11081 6620
rect 9751 5567 11081 5620
rect 11169 5567 11231 6673
rect 9751 5500 11231 5567
rect 11365 6673 12845 6740
rect 11365 6620 12695 6673
rect 11365 5620 11485 6620
rect 12485 5620 12695 6620
rect 11365 5567 12695 5620
rect 12783 5567 12845 6673
rect 11365 5500 12845 5567
rect 12979 6673 14459 6740
rect 12979 6620 14309 6673
rect 12979 5620 13099 6620
rect 14099 5620 14309 6620
rect 12979 5567 14309 5620
rect 14397 5567 14459 6673
rect 12979 5500 14459 5567
rect 14593 6673 16073 6740
rect 14593 6620 15923 6673
rect 14593 5620 14713 6620
rect 15713 5620 15923 6620
rect 14593 5567 15923 5620
rect 16011 5567 16073 6673
rect 14593 5500 16073 5567
rect 16207 6673 17687 6740
rect 16207 6620 17537 6673
rect 16207 5620 16327 6620
rect 17327 5620 17537 6620
rect 16207 5567 17537 5620
rect 17625 5567 17687 6673
rect 16207 5500 17687 5567
rect -17687 5313 -16207 5380
rect -17687 5260 -16357 5313
rect -17687 4260 -17567 5260
rect -16567 4260 -16357 5260
rect -17687 4207 -16357 4260
rect -16269 4207 -16207 5313
rect -17687 4140 -16207 4207
rect -16073 5313 -14593 5380
rect -16073 5260 -14743 5313
rect -16073 4260 -15953 5260
rect -14953 4260 -14743 5260
rect -16073 4207 -14743 4260
rect -14655 4207 -14593 5313
rect -16073 4140 -14593 4207
rect -14459 5313 -12979 5380
rect -14459 5260 -13129 5313
rect -14459 4260 -14339 5260
rect -13339 4260 -13129 5260
rect -14459 4207 -13129 4260
rect -13041 4207 -12979 5313
rect -14459 4140 -12979 4207
rect -12845 5313 -11365 5380
rect -12845 5260 -11515 5313
rect -12845 4260 -12725 5260
rect -11725 4260 -11515 5260
rect -12845 4207 -11515 4260
rect -11427 4207 -11365 5313
rect -12845 4140 -11365 4207
rect -11231 5313 -9751 5380
rect -11231 5260 -9901 5313
rect -11231 4260 -11111 5260
rect -10111 4260 -9901 5260
rect -11231 4207 -9901 4260
rect -9813 4207 -9751 5313
rect -11231 4140 -9751 4207
rect -9617 5313 -8137 5380
rect -9617 5260 -8287 5313
rect -9617 4260 -9497 5260
rect -8497 4260 -8287 5260
rect -9617 4207 -8287 4260
rect -8199 4207 -8137 5313
rect -9617 4140 -8137 4207
rect -8003 5313 -6523 5380
rect -8003 5260 -6673 5313
rect -8003 4260 -7883 5260
rect -6883 4260 -6673 5260
rect -8003 4207 -6673 4260
rect -6585 4207 -6523 5313
rect -8003 4140 -6523 4207
rect -6389 5313 -4909 5380
rect -6389 5260 -5059 5313
rect -6389 4260 -6269 5260
rect -5269 4260 -5059 5260
rect -6389 4207 -5059 4260
rect -4971 4207 -4909 5313
rect -6389 4140 -4909 4207
rect -4775 5313 -3295 5380
rect -4775 5260 -3445 5313
rect -4775 4260 -4655 5260
rect -3655 4260 -3445 5260
rect -4775 4207 -3445 4260
rect -3357 4207 -3295 5313
rect -4775 4140 -3295 4207
rect -3161 5313 -1681 5380
rect -3161 5260 -1831 5313
rect -3161 4260 -3041 5260
rect -2041 4260 -1831 5260
rect -3161 4207 -1831 4260
rect -1743 4207 -1681 5313
rect -3161 4140 -1681 4207
rect -1547 5313 -67 5380
rect -1547 5260 -217 5313
rect -1547 4260 -1427 5260
rect -427 4260 -217 5260
rect -1547 4207 -217 4260
rect -129 4207 -67 5313
rect -1547 4140 -67 4207
rect 67 5313 1547 5380
rect 67 5260 1397 5313
rect 67 4260 187 5260
rect 1187 4260 1397 5260
rect 67 4207 1397 4260
rect 1485 4207 1547 5313
rect 67 4140 1547 4207
rect 1681 5313 3161 5380
rect 1681 5260 3011 5313
rect 1681 4260 1801 5260
rect 2801 4260 3011 5260
rect 1681 4207 3011 4260
rect 3099 4207 3161 5313
rect 1681 4140 3161 4207
rect 3295 5313 4775 5380
rect 3295 5260 4625 5313
rect 3295 4260 3415 5260
rect 4415 4260 4625 5260
rect 3295 4207 4625 4260
rect 4713 4207 4775 5313
rect 3295 4140 4775 4207
rect 4909 5313 6389 5380
rect 4909 5260 6239 5313
rect 4909 4260 5029 5260
rect 6029 4260 6239 5260
rect 4909 4207 6239 4260
rect 6327 4207 6389 5313
rect 4909 4140 6389 4207
rect 6523 5313 8003 5380
rect 6523 5260 7853 5313
rect 6523 4260 6643 5260
rect 7643 4260 7853 5260
rect 6523 4207 7853 4260
rect 7941 4207 8003 5313
rect 6523 4140 8003 4207
rect 8137 5313 9617 5380
rect 8137 5260 9467 5313
rect 8137 4260 8257 5260
rect 9257 4260 9467 5260
rect 8137 4207 9467 4260
rect 9555 4207 9617 5313
rect 8137 4140 9617 4207
rect 9751 5313 11231 5380
rect 9751 5260 11081 5313
rect 9751 4260 9871 5260
rect 10871 4260 11081 5260
rect 9751 4207 11081 4260
rect 11169 4207 11231 5313
rect 9751 4140 11231 4207
rect 11365 5313 12845 5380
rect 11365 5260 12695 5313
rect 11365 4260 11485 5260
rect 12485 4260 12695 5260
rect 11365 4207 12695 4260
rect 12783 4207 12845 5313
rect 11365 4140 12845 4207
rect 12979 5313 14459 5380
rect 12979 5260 14309 5313
rect 12979 4260 13099 5260
rect 14099 4260 14309 5260
rect 12979 4207 14309 4260
rect 14397 4207 14459 5313
rect 12979 4140 14459 4207
rect 14593 5313 16073 5380
rect 14593 5260 15923 5313
rect 14593 4260 14713 5260
rect 15713 4260 15923 5260
rect 14593 4207 15923 4260
rect 16011 4207 16073 5313
rect 14593 4140 16073 4207
rect 16207 5313 17687 5380
rect 16207 5260 17537 5313
rect 16207 4260 16327 5260
rect 17327 4260 17537 5260
rect 16207 4207 17537 4260
rect 17625 4207 17687 5313
rect 16207 4140 17687 4207
rect -17687 3953 -16207 4020
rect -17687 3900 -16357 3953
rect -17687 2900 -17567 3900
rect -16567 2900 -16357 3900
rect -17687 2847 -16357 2900
rect -16269 2847 -16207 3953
rect -17687 2780 -16207 2847
rect -16073 3953 -14593 4020
rect -16073 3900 -14743 3953
rect -16073 2900 -15953 3900
rect -14953 2900 -14743 3900
rect -16073 2847 -14743 2900
rect -14655 2847 -14593 3953
rect -16073 2780 -14593 2847
rect -14459 3953 -12979 4020
rect -14459 3900 -13129 3953
rect -14459 2900 -14339 3900
rect -13339 2900 -13129 3900
rect -14459 2847 -13129 2900
rect -13041 2847 -12979 3953
rect -14459 2780 -12979 2847
rect -12845 3953 -11365 4020
rect -12845 3900 -11515 3953
rect -12845 2900 -12725 3900
rect -11725 2900 -11515 3900
rect -12845 2847 -11515 2900
rect -11427 2847 -11365 3953
rect -12845 2780 -11365 2847
rect -11231 3953 -9751 4020
rect -11231 3900 -9901 3953
rect -11231 2900 -11111 3900
rect -10111 2900 -9901 3900
rect -11231 2847 -9901 2900
rect -9813 2847 -9751 3953
rect -11231 2780 -9751 2847
rect -9617 3953 -8137 4020
rect -9617 3900 -8287 3953
rect -9617 2900 -9497 3900
rect -8497 2900 -8287 3900
rect -9617 2847 -8287 2900
rect -8199 2847 -8137 3953
rect -9617 2780 -8137 2847
rect -8003 3953 -6523 4020
rect -8003 3900 -6673 3953
rect -8003 2900 -7883 3900
rect -6883 2900 -6673 3900
rect -8003 2847 -6673 2900
rect -6585 2847 -6523 3953
rect -8003 2780 -6523 2847
rect -6389 3953 -4909 4020
rect -6389 3900 -5059 3953
rect -6389 2900 -6269 3900
rect -5269 2900 -5059 3900
rect -6389 2847 -5059 2900
rect -4971 2847 -4909 3953
rect -6389 2780 -4909 2847
rect -4775 3953 -3295 4020
rect -4775 3900 -3445 3953
rect -4775 2900 -4655 3900
rect -3655 2900 -3445 3900
rect -4775 2847 -3445 2900
rect -3357 2847 -3295 3953
rect -4775 2780 -3295 2847
rect -3161 3953 -1681 4020
rect -3161 3900 -1831 3953
rect -3161 2900 -3041 3900
rect -2041 2900 -1831 3900
rect -3161 2847 -1831 2900
rect -1743 2847 -1681 3953
rect -3161 2780 -1681 2847
rect -1547 3953 -67 4020
rect -1547 3900 -217 3953
rect -1547 2900 -1427 3900
rect -427 2900 -217 3900
rect -1547 2847 -217 2900
rect -129 2847 -67 3953
rect -1547 2780 -67 2847
rect 67 3953 1547 4020
rect 67 3900 1397 3953
rect 67 2900 187 3900
rect 1187 2900 1397 3900
rect 67 2847 1397 2900
rect 1485 2847 1547 3953
rect 67 2780 1547 2847
rect 1681 3953 3161 4020
rect 1681 3900 3011 3953
rect 1681 2900 1801 3900
rect 2801 2900 3011 3900
rect 1681 2847 3011 2900
rect 3099 2847 3161 3953
rect 1681 2780 3161 2847
rect 3295 3953 4775 4020
rect 3295 3900 4625 3953
rect 3295 2900 3415 3900
rect 4415 2900 4625 3900
rect 3295 2847 4625 2900
rect 4713 2847 4775 3953
rect 3295 2780 4775 2847
rect 4909 3953 6389 4020
rect 4909 3900 6239 3953
rect 4909 2900 5029 3900
rect 6029 2900 6239 3900
rect 4909 2847 6239 2900
rect 6327 2847 6389 3953
rect 4909 2780 6389 2847
rect 6523 3953 8003 4020
rect 6523 3900 7853 3953
rect 6523 2900 6643 3900
rect 7643 2900 7853 3900
rect 6523 2847 7853 2900
rect 7941 2847 8003 3953
rect 6523 2780 8003 2847
rect 8137 3953 9617 4020
rect 8137 3900 9467 3953
rect 8137 2900 8257 3900
rect 9257 2900 9467 3900
rect 8137 2847 9467 2900
rect 9555 2847 9617 3953
rect 8137 2780 9617 2847
rect 9751 3953 11231 4020
rect 9751 3900 11081 3953
rect 9751 2900 9871 3900
rect 10871 2900 11081 3900
rect 9751 2847 11081 2900
rect 11169 2847 11231 3953
rect 9751 2780 11231 2847
rect 11365 3953 12845 4020
rect 11365 3900 12695 3953
rect 11365 2900 11485 3900
rect 12485 2900 12695 3900
rect 11365 2847 12695 2900
rect 12783 2847 12845 3953
rect 11365 2780 12845 2847
rect 12979 3953 14459 4020
rect 12979 3900 14309 3953
rect 12979 2900 13099 3900
rect 14099 2900 14309 3900
rect 12979 2847 14309 2900
rect 14397 2847 14459 3953
rect 12979 2780 14459 2847
rect 14593 3953 16073 4020
rect 14593 3900 15923 3953
rect 14593 2900 14713 3900
rect 15713 2900 15923 3900
rect 14593 2847 15923 2900
rect 16011 2847 16073 3953
rect 14593 2780 16073 2847
rect 16207 3953 17687 4020
rect 16207 3900 17537 3953
rect 16207 2900 16327 3900
rect 17327 2900 17537 3900
rect 16207 2847 17537 2900
rect 17625 2847 17687 3953
rect 16207 2780 17687 2847
rect -17687 2593 -16207 2660
rect -17687 2540 -16357 2593
rect -17687 1540 -17567 2540
rect -16567 1540 -16357 2540
rect -17687 1487 -16357 1540
rect -16269 1487 -16207 2593
rect -17687 1420 -16207 1487
rect -16073 2593 -14593 2660
rect -16073 2540 -14743 2593
rect -16073 1540 -15953 2540
rect -14953 1540 -14743 2540
rect -16073 1487 -14743 1540
rect -14655 1487 -14593 2593
rect -16073 1420 -14593 1487
rect -14459 2593 -12979 2660
rect -14459 2540 -13129 2593
rect -14459 1540 -14339 2540
rect -13339 1540 -13129 2540
rect -14459 1487 -13129 1540
rect -13041 1487 -12979 2593
rect -14459 1420 -12979 1487
rect -12845 2593 -11365 2660
rect -12845 2540 -11515 2593
rect -12845 1540 -12725 2540
rect -11725 1540 -11515 2540
rect -12845 1487 -11515 1540
rect -11427 1487 -11365 2593
rect -12845 1420 -11365 1487
rect -11231 2593 -9751 2660
rect -11231 2540 -9901 2593
rect -11231 1540 -11111 2540
rect -10111 1540 -9901 2540
rect -11231 1487 -9901 1540
rect -9813 1487 -9751 2593
rect -11231 1420 -9751 1487
rect -9617 2593 -8137 2660
rect -9617 2540 -8287 2593
rect -9617 1540 -9497 2540
rect -8497 1540 -8287 2540
rect -9617 1487 -8287 1540
rect -8199 1487 -8137 2593
rect -9617 1420 -8137 1487
rect -8003 2593 -6523 2660
rect -8003 2540 -6673 2593
rect -8003 1540 -7883 2540
rect -6883 1540 -6673 2540
rect -8003 1487 -6673 1540
rect -6585 1487 -6523 2593
rect -8003 1420 -6523 1487
rect -6389 2593 -4909 2660
rect -6389 2540 -5059 2593
rect -6389 1540 -6269 2540
rect -5269 1540 -5059 2540
rect -6389 1487 -5059 1540
rect -4971 1487 -4909 2593
rect -6389 1420 -4909 1487
rect -4775 2593 -3295 2660
rect -4775 2540 -3445 2593
rect -4775 1540 -4655 2540
rect -3655 1540 -3445 2540
rect -4775 1487 -3445 1540
rect -3357 1487 -3295 2593
rect -4775 1420 -3295 1487
rect -3161 2593 -1681 2660
rect -3161 2540 -1831 2593
rect -3161 1540 -3041 2540
rect -2041 1540 -1831 2540
rect -3161 1487 -1831 1540
rect -1743 1487 -1681 2593
rect -3161 1420 -1681 1487
rect -1547 2593 -67 2660
rect -1547 2540 -217 2593
rect -1547 1540 -1427 2540
rect -427 1540 -217 2540
rect -1547 1487 -217 1540
rect -129 1487 -67 2593
rect -1547 1420 -67 1487
rect 67 2593 1547 2660
rect 67 2540 1397 2593
rect 67 1540 187 2540
rect 1187 1540 1397 2540
rect 67 1487 1397 1540
rect 1485 1487 1547 2593
rect 67 1420 1547 1487
rect 1681 2593 3161 2660
rect 1681 2540 3011 2593
rect 1681 1540 1801 2540
rect 2801 1540 3011 2540
rect 1681 1487 3011 1540
rect 3099 1487 3161 2593
rect 1681 1420 3161 1487
rect 3295 2593 4775 2660
rect 3295 2540 4625 2593
rect 3295 1540 3415 2540
rect 4415 1540 4625 2540
rect 3295 1487 4625 1540
rect 4713 1487 4775 2593
rect 3295 1420 4775 1487
rect 4909 2593 6389 2660
rect 4909 2540 6239 2593
rect 4909 1540 5029 2540
rect 6029 1540 6239 2540
rect 4909 1487 6239 1540
rect 6327 1487 6389 2593
rect 4909 1420 6389 1487
rect 6523 2593 8003 2660
rect 6523 2540 7853 2593
rect 6523 1540 6643 2540
rect 7643 1540 7853 2540
rect 6523 1487 7853 1540
rect 7941 1487 8003 2593
rect 6523 1420 8003 1487
rect 8137 2593 9617 2660
rect 8137 2540 9467 2593
rect 8137 1540 8257 2540
rect 9257 1540 9467 2540
rect 8137 1487 9467 1540
rect 9555 1487 9617 2593
rect 8137 1420 9617 1487
rect 9751 2593 11231 2660
rect 9751 2540 11081 2593
rect 9751 1540 9871 2540
rect 10871 1540 11081 2540
rect 9751 1487 11081 1540
rect 11169 1487 11231 2593
rect 9751 1420 11231 1487
rect 11365 2593 12845 2660
rect 11365 2540 12695 2593
rect 11365 1540 11485 2540
rect 12485 1540 12695 2540
rect 11365 1487 12695 1540
rect 12783 1487 12845 2593
rect 11365 1420 12845 1487
rect 12979 2593 14459 2660
rect 12979 2540 14309 2593
rect 12979 1540 13099 2540
rect 14099 1540 14309 2540
rect 12979 1487 14309 1540
rect 14397 1487 14459 2593
rect 12979 1420 14459 1487
rect 14593 2593 16073 2660
rect 14593 2540 15923 2593
rect 14593 1540 14713 2540
rect 15713 1540 15923 2540
rect 14593 1487 15923 1540
rect 16011 1487 16073 2593
rect 14593 1420 16073 1487
rect 16207 2593 17687 2660
rect 16207 2540 17537 2593
rect 16207 1540 16327 2540
rect 17327 1540 17537 2540
rect 16207 1487 17537 1540
rect 17625 1487 17687 2593
rect 16207 1420 17687 1487
rect -17687 1233 -16207 1300
rect -17687 1180 -16357 1233
rect -17687 180 -17567 1180
rect -16567 180 -16357 1180
rect -17687 127 -16357 180
rect -16269 127 -16207 1233
rect -17687 60 -16207 127
rect -16073 1233 -14593 1300
rect -16073 1180 -14743 1233
rect -16073 180 -15953 1180
rect -14953 180 -14743 1180
rect -16073 127 -14743 180
rect -14655 127 -14593 1233
rect -16073 60 -14593 127
rect -14459 1233 -12979 1300
rect -14459 1180 -13129 1233
rect -14459 180 -14339 1180
rect -13339 180 -13129 1180
rect -14459 127 -13129 180
rect -13041 127 -12979 1233
rect -14459 60 -12979 127
rect -12845 1233 -11365 1300
rect -12845 1180 -11515 1233
rect -12845 180 -12725 1180
rect -11725 180 -11515 1180
rect -12845 127 -11515 180
rect -11427 127 -11365 1233
rect -12845 60 -11365 127
rect -11231 1233 -9751 1300
rect -11231 1180 -9901 1233
rect -11231 180 -11111 1180
rect -10111 180 -9901 1180
rect -11231 127 -9901 180
rect -9813 127 -9751 1233
rect -11231 60 -9751 127
rect -9617 1233 -8137 1300
rect -9617 1180 -8287 1233
rect -9617 180 -9497 1180
rect -8497 180 -8287 1180
rect -9617 127 -8287 180
rect -8199 127 -8137 1233
rect -9617 60 -8137 127
rect -8003 1233 -6523 1300
rect -8003 1180 -6673 1233
rect -8003 180 -7883 1180
rect -6883 180 -6673 1180
rect -8003 127 -6673 180
rect -6585 127 -6523 1233
rect -8003 60 -6523 127
rect -6389 1233 -4909 1300
rect -6389 1180 -5059 1233
rect -6389 180 -6269 1180
rect -5269 180 -5059 1180
rect -6389 127 -5059 180
rect -4971 127 -4909 1233
rect -6389 60 -4909 127
rect -4775 1233 -3295 1300
rect -4775 1180 -3445 1233
rect -4775 180 -4655 1180
rect -3655 180 -3445 1180
rect -4775 127 -3445 180
rect -3357 127 -3295 1233
rect -4775 60 -3295 127
rect -3161 1233 -1681 1300
rect -3161 1180 -1831 1233
rect -3161 180 -3041 1180
rect -2041 180 -1831 1180
rect -3161 127 -1831 180
rect -1743 127 -1681 1233
rect -3161 60 -1681 127
rect -1547 1233 -67 1300
rect -1547 1180 -217 1233
rect -1547 180 -1427 1180
rect -427 180 -217 1180
rect -1547 127 -217 180
rect -129 127 -67 1233
rect -1547 60 -67 127
rect 67 1233 1547 1300
rect 67 1180 1397 1233
rect 67 180 187 1180
rect 1187 180 1397 1180
rect 67 127 1397 180
rect 1485 127 1547 1233
rect 67 60 1547 127
rect 1681 1233 3161 1300
rect 1681 1180 3011 1233
rect 1681 180 1801 1180
rect 2801 180 3011 1180
rect 1681 127 3011 180
rect 3099 127 3161 1233
rect 1681 60 3161 127
rect 3295 1233 4775 1300
rect 3295 1180 4625 1233
rect 3295 180 3415 1180
rect 4415 180 4625 1180
rect 3295 127 4625 180
rect 4713 127 4775 1233
rect 3295 60 4775 127
rect 4909 1233 6389 1300
rect 4909 1180 6239 1233
rect 4909 180 5029 1180
rect 6029 180 6239 1180
rect 4909 127 6239 180
rect 6327 127 6389 1233
rect 4909 60 6389 127
rect 6523 1233 8003 1300
rect 6523 1180 7853 1233
rect 6523 180 6643 1180
rect 7643 180 7853 1180
rect 6523 127 7853 180
rect 7941 127 8003 1233
rect 6523 60 8003 127
rect 8137 1233 9617 1300
rect 8137 1180 9467 1233
rect 8137 180 8257 1180
rect 9257 180 9467 1180
rect 8137 127 9467 180
rect 9555 127 9617 1233
rect 8137 60 9617 127
rect 9751 1233 11231 1300
rect 9751 1180 11081 1233
rect 9751 180 9871 1180
rect 10871 180 11081 1180
rect 9751 127 11081 180
rect 11169 127 11231 1233
rect 9751 60 11231 127
rect 11365 1233 12845 1300
rect 11365 1180 12695 1233
rect 11365 180 11485 1180
rect 12485 180 12695 1180
rect 11365 127 12695 180
rect 12783 127 12845 1233
rect 11365 60 12845 127
rect 12979 1233 14459 1300
rect 12979 1180 14309 1233
rect 12979 180 13099 1180
rect 14099 180 14309 1180
rect 12979 127 14309 180
rect 14397 127 14459 1233
rect 12979 60 14459 127
rect 14593 1233 16073 1300
rect 14593 1180 15923 1233
rect 14593 180 14713 1180
rect 15713 180 15923 1180
rect 14593 127 15923 180
rect 16011 127 16073 1233
rect 14593 60 16073 127
rect 16207 1233 17687 1300
rect 16207 1180 17537 1233
rect 16207 180 16327 1180
rect 17327 180 17537 1180
rect 16207 127 17537 180
rect 17625 127 17687 1233
rect 16207 60 17687 127
rect -17687 -127 -16207 -60
rect -17687 -180 -16357 -127
rect -17687 -1180 -17567 -180
rect -16567 -1180 -16357 -180
rect -17687 -1233 -16357 -1180
rect -16269 -1233 -16207 -127
rect -17687 -1300 -16207 -1233
rect -16073 -127 -14593 -60
rect -16073 -180 -14743 -127
rect -16073 -1180 -15953 -180
rect -14953 -1180 -14743 -180
rect -16073 -1233 -14743 -1180
rect -14655 -1233 -14593 -127
rect -16073 -1300 -14593 -1233
rect -14459 -127 -12979 -60
rect -14459 -180 -13129 -127
rect -14459 -1180 -14339 -180
rect -13339 -1180 -13129 -180
rect -14459 -1233 -13129 -1180
rect -13041 -1233 -12979 -127
rect -14459 -1300 -12979 -1233
rect -12845 -127 -11365 -60
rect -12845 -180 -11515 -127
rect -12845 -1180 -12725 -180
rect -11725 -1180 -11515 -180
rect -12845 -1233 -11515 -1180
rect -11427 -1233 -11365 -127
rect -12845 -1300 -11365 -1233
rect -11231 -127 -9751 -60
rect -11231 -180 -9901 -127
rect -11231 -1180 -11111 -180
rect -10111 -1180 -9901 -180
rect -11231 -1233 -9901 -1180
rect -9813 -1233 -9751 -127
rect -11231 -1300 -9751 -1233
rect -9617 -127 -8137 -60
rect -9617 -180 -8287 -127
rect -9617 -1180 -9497 -180
rect -8497 -1180 -8287 -180
rect -9617 -1233 -8287 -1180
rect -8199 -1233 -8137 -127
rect -9617 -1300 -8137 -1233
rect -8003 -127 -6523 -60
rect -8003 -180 -6673 -127
rect -8003 -1180 -7883 -180
rect -6883 -1180 -6673 -180
rect -8003 -1233 -6673 -1180
rect -6585 -1233 -6523 -127
rect -8003 -1300 -6523 -1233
rect -6389 -127 -4909 -60
rect -6389 -180 -5059 -127
rect -6389 -1180 -6269 -180
rect -5269 -1180 -5059 -180
rect -6389 -1233 -5059 -1180
rect -4971 -1233 -4909 -127
rect -6389 -1300 -4909 -1233
rect -4775 -127 -3295 -60
rect -4775 -180 -3445 -127
rect -4775 -1180 -4655 -180
rect -3655 -1180 -3445 -180
rect -4775 -1233 -3445 -1180
rect -3357 -1233 -3295 -127
rect -4775 -1300 -3295 -1233
rect -3161 -127 -1681 -60
rect -3161 -180 -1831 -127
rect -3161 -1180 -3041 -180
rect -2041 -1180 -1831 -180
rect -3161 -1233 -1831 -1180
rect -1743 -1233 -1681 -127
rect -3161 -1300 -1681 -1233
rect -1547 -127 -67 -60
rect -1547 -180 -217 -127
rect -1547 -1180 -1427 -180
rect -427 -1180 -217 -180
rect -1547 -1233 -217 -1180
rect -129 -1233 -67 -127
rect -1547 -1300 -67 -1233
rect 67 -127 1547 -60
rect 67 -180 1397 -127
rect 67 -1180 187 -180
rect 1187 -1180 1397 -180
rect 67 -1233 1397 -1180
rect 1485 -1233 1547 -127
rect 67 -1300 1547 -1233
rect 1681 -127 3161 -60
rect 1681 -180 3011 -127
rect 1681 -1180 1801 -180
rect 2801 -1180 3011 -180
rect 1681 -1233 3011 -1180
rect 3099 -1233 3161 -127
rect 1681 -1300 3161 -1233
rect 3295 -127 4775 -60
rect 3295 -180 4625 -127
rect 3295 -1180 3415 -180
rect 4415 -1180 4625 -180
rect 3295 -1233 4625 -1180
rect 4713 -1233 4775 -127
rect 3295 -1300 4775 -1233
rect 4909 -127 6389 -60
rect 4909 -180 6239 -127
rect 4909 -1180 5029 -180
rect 6029 -1180 6239 -180
rect 4909 -1233 6239 -1180
rect 6327 -1233 6389 -127
rect 4909 -1300 6389 -1233
rect 6523 -127 8003 -60
rect 6523 -180 7853 -127
rect 6523 -1180 6643 -180
rect 7643 -1180 7853 -180
rect 6523 -1233 7853 -1180
rect 7941 -1233 8003 -127
rect 6523 -1300 8003 -1233
rect 8137 -127 9617 -60
rect 8137 -180 9467 -127
rect 8137 -1180 8257 -180
rect 9257 -1180 9467 -180
rect 8137 -1233 9467 -1180
rect 9555 -1233 9617 -127
rect 8137 -1300 9617 -1233
rect 9751 -127 11231 -60
rect 9751 -180 11081 -127
rect 9751 -1180 9871 -180
rect 10871 -1180 11081 -180
rect 9751 -1233 11081 -1180
rect 11169 -1233 11231 -127
rect 9751 -1300 11231 -1233
rect 11365 -127 12845 -60
rect 11365 -180 12695 -127
rect 11365 -1180 11485 -180
rect 12485 -1180 12695 -180
rect 11365 -1233 12695 -1180
rect 12783 -1233 12845 -127
rect 11365 -1300 12845 -1233
rect 12979 -127 14459 -60
rect 12979 -180 14309 -127
rect 12979 -1180 13099 -180
rect 14099 -1180 14309 -180
rect 12979 -1233 14309 -1180
rect 14397 -1233 14459 -127
rect 12979 -1300 14459 -1233
rect 14593 -127 16073 -60
rect 14593 -180 15923 -127
rect 14593 -1180 14713 -180
rect 15713 -1180 15923 -180
rect 14593 -1233 15923 -1180
rect 16011 -1233 16073 -127
rect 14593 -1300 16073 -1233
rect 16207 -127 17687 -60
rect 16207 -180 17537 -127
rect 16207 -1180 16327 -180
rect 17327 -1180 17537 -180
rect 16207 -1233 17537 -1180
rect 17625 -1233 17687 -127
rect 16207 -1300 17687 -1233
rect -17687 -1487 -16207 -1420
rect -17687 -1540 -16357 -1487
rect -17687 -2540 -17567 -1540
rect -16567 -2540 -16357 -1540
rect -17687 -2593 -16357 -2540
rect -16269 -2593 -16207 -1487
rect -17687 -2660 -16207 -2593
rect -16073 -1487 -14593 -1420
rect -16073 -1540 -14743 -1487
rect -16073 -2540 -15953 -1540
rect -14953 -2540 -14743 -1540
rect -16073 -2593 -14743 -2540
rect -14655 -2593 -14593 -1487
rect -16073 -2660 -14593 -2593
rect -14459 -1487 -12979 -1420
rect -14459 -1540 -13129 -1487
rect -14459 -2540 -14339 -1540
rect -13339 -2540 -13129 -1540
rect -14459 -2593 -13129 -2540
rect -13041 -2593 -12979 -1487
rect -14459 -2660 -12979 -2593
rect -12845 -1487 -11365 -1420
rect -12845 -1540 -11515 -1487
rect -12845 -2540 -12725 -1540
rect -11725 -2540 -11515 -1540
rect -12845 -2593 -11515 -2540
rect -11427 -2593 -11365 -1487
rect -12845 -2660 -11365 -2593
rect -11231 -1487 -9751 -1420
rect -11231 -1540 -9901 -1487
rect -11231 -2540 -11111 -1540
rect -10111 -2540 -9901 -1540
rect -11231 -2593 -9901 -2540
rect -9813 -2593 -9751 -1487
rect -11231 -2660 -9751 -2593
rect -9617 -1487 -8137 -1420
rect -9617 -1540 -8287 -1487
rect -9617 -2540 -9497 -1540
rect -8497 -2540 -8287 -1540
rect -9617 -2593 -8287 -2540
rect -8199 -2593 -8137 -1487
rect -9617 -2660 -8137 -2593
rect -8003 -1487 -6523 -1420
rect -8003 -1540 -6673 -1487
rect -8003 -2540 -7883 -1540
rect -6883 -2540 -6673 -1540
rect -8003 -2593 -6673 -2540
rect -6585 -2593 -6523 -1487
rect -8003 -2660 -6523 -2593
rect -6389 -1487 -4909 -1420
rect -6389 -1540 -5059 -1487
rect -6389 -2540 -6269 -1540
rect -5269 -2540 -5059 -1540
rect -6389 -2593 -5059 -2540
rect -4971 -2593 -4909 -1487
rect -6389 -2660 -4909 -2593
rect -4775 -1487 -3295 -1420
rect -4775 -1540 -3445 -1487
rect -4775 -2540 -4655 -1540
rect -3655 -2540 -3445 -1540
rect -4775 -2593 -3445 -2540
rect -3357 -2593 -3295 -1487
rect -4775 -2660 -3295 -2593
rect -3161 -1487 -1681 -1420
rect -3161 -1540 -1831 -1487
rect -3161 -2540 -3041 -1540
rect -2041 -2540 -1831 -1540
rect -3161 -2593 -1831 -2540
rect -1743 -2593 -1681 -1487
rect -3161 -2660 -1681 -2593
rect -1547 -1487 -67 -1420
rect -1547 -1540 -217 -1487
rect -1547 -2540 -1427 -1540
rect -427 -2540 -217 -1540
rect -1547 -2593 -217 -2540
rect -129 -2593 -67 -1487
rect -1547 -2660 -67 -2593
rect 67 -1487 1547 -1420
rect 67 -1540 1397 -1487
rect 67 -2540 187 -1540
rect 1187 -2540 1397 -1540
rect 67 -2593 1397 -2540
rect 1485 -2593 1547 -1487
rect 67 -2660 1547 -2593
rect 1681 -1487 3161 -1420
rect 1681 -1540 3011 -1487
rect 1681 -2540 1801 -1540
rect 2801 -2540 3011 -1540
rect 1681 -2593 3011 -2540
rect 3099 -2593 3161 -1487
rect 1681 -2660 3161 -2593
rect 3295 -1487 4775 -1420
rect 3295 -1540 4625 -1487
rect 3295 -2540 3415 -1540
rect 4415 -2540 4625 -1540
rect 3295 -2593 4625 -2540
rect 4713 -2593 4775 -1487
rect 3295 -2660 4775 -2593
rect 4909 -1487 6389 -1420
rect 4909 -1540 6239 -1487
rect 4909 -2540 5029 -1540
rect 6029 -2540 6239 -1540
rect 4909 -2593 6239 -2540
rect 6327 -2593 6389 -1487
rect 4909 -2660 6389 -2593
rect 6523 -1487 8003 -1420
rect 6523 -1540 7853 -1487
rect 6523 -2540 6643 -1540
rect 7643 -2540 7853 -1540
rect 6523 -2593 7853 -2540
rect 7941 -2593 8003 -1487
rect 6523 -2660 8003 -2593
rect 8137 -1487 9617 -1420
rect 8137 -1540 9467 -1487
rect 8137 -2540 8257 -1540
rect 9257 -2540 9467 -1540
rect 8137 -2593 9467 -2540
rect 9555 -2593 9617 -1487
rect 8137 -2660 9617 -2593
rect 9751 -1487 11231 -1420
rect 9751 -1540 11081 -1487
rect 9751 -2540 9871 -1540
rect 10871 -2540 11081 -1540
rect 9751 -2593 11081 -2540
rect 11169 -2593 11231 -1487
rect 9751 -2660 11231 -2593
rect 11365 -1487 12845 -1420
rect 11365 -1540 12695 -1487
rect 11365 -2540 11485 -1540
rect 12485 -2540 12695 -1540
rect 11365 -2593 12695 -2540
rect 12783 -2593 12845 -1487
rect 11365 -2660 12845 -2593
rect 12979 -1487 14459 -1420
rect 12979 -1540 14309 -1487
rect 12979 -2540 13099 -1540
rect 14099 -2540 14309 -1540
rect 12979 -2593 14309 -2540
rect 14397 -2593 14459 -1487
rect 12979 -2660 14459 -2593
rect 14593 -1487 16073 -1420
rect 14593 -1540 15923 -1487
rect 14593 -2540 14713 -1540
rect 15713 -2540 15923 -1540
rect 14593 -2593 15923 -2540
rect 16011 -2593 16073 -1487
rect 14593 -2660 16073 -2593
rect 16207 -1487 17687 -1420
rect 16207 -1540 17537 -1487
rect 16207 -2540 16327 -1540
rect 17327 -2540 17537 -1540
rect 16207 -2593 17537 -2540
rect 17625 -2593 17687 -1487
rect 16207 -2660 17687 -2593
rect -17687 -2847 -16207 -2780
rect -17687 -2900 -16357 -2847
rect -17687 -3900 -17567 -2900
rect -16567 -3900 -16357 -2900
rect -17687 -3953 -16357 -3900
rect -16269 -3953 -16207 -2847
rect -17687 -4020 -16207 -3953
rect -16073 -2847 -14593 -2780
rect -16073 -2900 -14743 -2847
rect -16073 -3900 -15953 -2900
rect -14953 -3900 -14743 -2900
rect -16073 -3953 -14743 -3900
rect -14655 -3953 -14593 -2847
rect -16073 -4020 -14593 -3953
rect -14459 -2847 -12979 -2780
rect -14459 -2900 -13129 -2847
rect -14459 -3900 -14339 -2900
rect -13339 -3900 -13129 -2900
rect -14459 -3953 -13129 -3900
rect -13041 -3953 -12979 -2847
rect -14459 -4020 -12979 -3953
rect -12845 -2847 -11365 -2780
rect -12845 -2900 -11515 -2847
rect -12845 -3900 -12725 -2900
rect -11725 -3900 -11515 -2900
rect -12845 -3953 -11515 -3900
rect -11427 -3953 -11365 -2847
rect -12845 -4020 -11365 -3953
rect -11231 -2847 -9751 -2780
rect -11231 -2900 -9901 -2847
rect -11231 -3900 -11111 -2900
rect -10111 -3900 -9901 -2900
rect -11231 -3953 -9901 -3900
rect -9813 -3953 -9751 -2847
rect -11231 -4020 -9751 -3953
rect -9617 -2847 -8137 -2780
rect -9617 -2900 -8287 -2847
rect -9617 -3900 -9497 -2900
rect -8497 -3900 -8287 -2900
rect -9617 -3953 -8287 -3900
rect -8199 -3953 -8137 -2847
rect -9617 -4020 -8137 -3953
rect -8003 -2847 -6523 -2780
rect -8003 -2900 -6673 -2847
rect -8003 -3900 -7883 -2900
rect -6883 -3900 -6673 -2900
rect -8003 -3953 -6673 -3900
rect -6585 -3953 -6523 -2847
rect -8003 -4020 -6523 -3953
rect -6389 -2847 -4909 -2780
rect -6389 -2900 -5059 -2847
rect -6389 -3900 -6269 -2900
rect -5269 -3900 -5059 -2900
rect -6389 -3953 -5059 -3900
rect -4971 -3953 -4909 -2847
rect -6389 -4020 -4909 -3953
rect -4775 -2847 -3295 -2780
rect -4775 -2900 -3445 -2847
rect -4775 -3900 -4655 -2900
rect -3655 -3900 -3445 -2900
rect -4775 -3953 -3445 -3900
rect -3357 -3953 -3295 -2847
rect -4775 -4020 -3295 -3953
rect -3161 -2847 -1681 -2780
rect -3161 -2900 -1831 -2847
rect -3161 -3900 -3041 -2900
rect -2041 -3900 -1831 -2900
rect -3161 -3953 -1831 -3900
rect -1743 -3953 -1681 -2847
rect -3161 -4020 -1681 -3953
rect -1547 -2847 -67 -2780
rect -1547 -2900 -217 -2847
rect -1547 -3900 -1427 -2900
rect -427 -3900 -217 -2900
rect -1547 -3953 -217 -3900
rect -129 -3953 -67 -2847
rect -1547 -4020 -67 -3953
rect 67 -2847 1547 -2780
rect 67 -2900 1397 -2847
rect 67 -3900 187 -2900
rect 1187 -3900 1397 -2900
rect 67 -3953 1397 -3900
rect 1485 -3953 1547 -2847
rect 67 -4020 1547 -3953
rect 1681 -2847 3161 -2780
rect 1681 -2900 3011 -2847
rect 1681 -3900 1801 -2900
rect 2801 -3900 3011 -2900
rect 1681 -3953 3011 -3900
rect 3099 -3953 3161 -2847
rect 1681 -4020 3161 -3953
rect 3295 -2847 4775 -2780
rect 3295 -2900 4625 -2847
rect 3295 -3900 3415 -2900
rect 4415 -3900 4625 -2900
rect 3295 -3953 4625 -3900
rect 4713 -3953 4775 -2847
rect 3295 -4020 4775 -3953
rect 4909 -2847 6389 -2780
rect 4909 -2900 6239 -2847
rect 4909 -3900 5029 -2900
rect 6029 -3900 6239 -2900
rect 4909 -3953 6239 -3900
rect 6327 -3953 6389 -2847
rect 4909 -4020 6389 -3953
rect 6523 -2847 8003 -2780
rect 6523 -2900 7853 -2847
rect 6523 -3900 6643 -2900
rect 7643 -3900 7853 -2900
rect 6523 -3953 7853 -3900
rect 7941 -3953 8003 -2847
rect 6523 -4020 8003 -3953
rect 8137 -2847 9617 -2780
rect 8137 -2900 9467 -2847
rect 8137 -3900 8257 -2900
rect 9257 -3900 9467 -2900
rect 8137 -3953 9467 -3900
rect 9555 -3953 9617 -2847
rect 8137 -4020 9617 -3953
rect 9751 -2847 11231 -2780
rect 9751 -2900 11081 -2847
rect 9751 -3900 9871 -2900
rect 10871 -3900 11081 -2900
rect 9751 -3953 11081 -3900
rect 11169 -3953 11231 -2847
rect 9751 -4020 11231 -3953
rect 11365 -2847 12845 -2780
rect 11365 -2900 12695 -2847
rect 11365 -3900 11485 -2900
rect 12485 -3900 12695 -2900
rect 11365 -3953 12695 -3900
rect 12783 -3953 12845 -2847
rect 11365 -4020 12845 -3953
rect 12979 -2847 14459 -2780
rect 12979 -2900 14309 -2847
rect 12979 -3900 13099 -2900
rect 14099 -3900 14309 -2900
rect 12979 -3953 14309 -3900
rect 14397 -3953 14459 -2847
rect 12979 -4020 14459 -3953
rect 14593 -2847 16073 -2780
rect 14593 -2900 15923 -2847
rect 14593 -3900 14713 -2900
rect 15713 -3900 15923 -2900
rect 14593 -3953 15923 -3900
rect 16011 -3953 16073 -2847
rect 14593 -4020 16073 -3953
rect 16207 -2847 17687 -2780
rect 16207 -2900 17537 -2847
rect 16207 -3900 16327 -2900
rect 17327 -3900 17537 -2900
rect 16207 -3953 17537 -3900
rect 17625 -3953 17687 -2847
rect 16207 -4020 17687 -3953
rect -17687 -4207 -16207 -4140
rect -17687 -4260 -16357 -4207
rect -17687 -5260 -17567 -4260
rect -16567 -5260 -16357 -4260
rect -17687 -5313 -16357 -5260
rect -16269 -5313 -16207 -4207
rect -17687 -5380 -16207 -5313
rect -16073 -4207 -14593 -4140
rect -16073 -4260 -14743 -4207
rect -16073 -5260 -15953 -4260
rect -14953 -5260 -14743 -4260
rect -16073 -5313 -14743 -5260
rect -14655 -5313 -14593 -4207
rect -16073 -5380 -14593 -5313
rect -14459 -4207 -12979 -4140
rect -14459 -4260 -13129 -4207
rect -14459 -5260 -14339 -4260
rect -13339 -5260 -13129 -4260
rect -14459 -5313 -13129 -5260
rect -13041 -5313 -12979 -4207
rect -14459 -5380 -12979 -5313
rect -12845 -4207 -11365 -4140
rect -12845 -4260 -11515 -4207
rect -12845 -5260 -12725 -4260
rect -11725 -5260 -11515 -4260
rect -12845 -5313 -11515 -5260
rect -11427 -5313 -11365 -4207
rect -12845 -5380 -11365 -5313
rect -11231 -4207 -9751 -4140
rect -11231 -4260 -9901 -4207
rect -11231 -5260 -11111 -4260
rect -10111 -5260 -9901 -4260
rect -11231 -5313 -9901 -5260
rect -9813 -5313 -9751 -4207
rect -11231 -5380 -9751 -5313
rect -9617 -4207 -8137 -4140
rect -9617 -4260 -8287 -4207
rect -9617 -5260 -9497 -4260
rect -8497 -5260 -8287 -4260
rect -9617 -5313 -8287 -5260
rect -8199 -5313 -8137 -4207
rect -9617 -5380 -8137 -5313
rect -8003 -4207 -6523 -4140
rect -8003 -4260 -6673 -4207
rect -8003 -5260 -7883 -4260
rect -6883 -5260 -6673 -4260
rect -8003 -5313 -6673 -5260
rect -6585 -5313 -6523 -4207
rect -8003 -5380 -6523 -5313
rect -6389 -4207 -4909 -4140
rect -6389 -4260 -5059 -4207
rect -6389 -5260 -6269 -4260
rect -5269 -5260 -5059 -4260
rect -6389 -5313 -5059 -5260
rect -4971 -5313 -4909 -4207
rect -6389 -5380 -4909 -5313
rect -4775 -4207 -3295 -4140
rect -4775 -4260 -3445 -4207
rect -4775 -5260 -4655 -4260
rect -3655 -5260 -3445 -4260
rect -4775 -5313 -3445 -5260
rect -3357 -5313 -3295 -4207
rect -4775 -5380 -3295 -5313
rect -3161 -4207 -1681 -4140
rect -3161 -4260 -1831 -4207
rect -3161 -5260 -3041 -4260
rect -2041 -5260 -1831 -4260
rect -3161 -5313 -1831 -5260
rect -1743 -5313 -1681 -4207
rect -3161 -5380 -1681 -5313
rect -1547 -4207 -67 -4140
rect -1547 -4260 -217 -4207
rect -1547 -5260 -1427 -4260
rect -427 -5260 -217 -4260
rect -1547 -5313 -217 -5260
rect -129 -5313 -67 -4207
rect -1547 -5380 -67 -5313
rect 67 -4207 1547 -4140
rect 67 -4260 1397 -4207
rect 67 -5260 187 -4260
rect 1187 -5260 1397 -4260
rect 67 -5313 1397 -5260
rect 1485 -5313 1547 -4207
rect 67 -5380 1547 -5313
rect 1681 -4207 3161 -4140
rect 1681 -4260 3011 -4207
rect 1681 -5260 1801 -4260
rect 2801 -5260 3011 -4260
rect 1681 -5313 3011 -5260
rect 3099 -5313 3161 -4207
rect 1681 -5380 3161 -5313
rect 3295 -4207 4775 -4140
rect 3295 -4260 4625 -4207
rect 3295 -5260 3415 -4260
rect 4415 -5260 4625 -4260
rect 3295 -5313 4625 -5260
rect 4713 -5313 4775 -4207
rect 3295 -5380 4775 -5313
rect 4909 -4207 6389 -4140
rect 4909 -4260 6239 -4207
rect 4909 -5260 5029 -4260
rect 6029 -5260 6239 -4260
rect 4909 -5313 6239 -5260
rect 6327 -5313 6389 -4207
rect 4909 -5380 6389 -5313
rect 6523 -4207 8003 -4140
rect 6523 -4260 7853 -4207
rect 6523 -5260 6643 -4260
rect 7643 -5260 7853 -4260
rect 6523 -5313 7853 -5260
rect 7941 -5313 8003 -4207
rect 6523 -5380 8003 -5313
rect 8137 -4207 9617 -4140
rect 8137 -4260 9467 -4207
rect 8137 -5260 8257 -4260
rect 9257 -5260 9467 -4260
rect 8137 -5313 9467 -5260
rect 9555 -5313 9617 -4207
rect 8137 -5380 9617 -5313
rect 9751 -4207 11231 -4140
rect 9751 -4260 11081 -4207
rect 9751 -5260 9871 -4260
rect 10871 -5260 11081 -4260
rect 9751 -5313 11081 -5260
rect 11169 -5313 11231 -4207
rect 9751 -5380 11231 -5313
rect 11365 -4207 12845 -4140
rect 11365 -4260 12695 -4207
rect 11365 -5260 11485 -4260
rect 12485 -5260 12695 -4260
rect 11365 -5313 12695 -5260
rect 12783 -5313 12845 -4207
rect 11365 -5380 12845 -5313
rect 12979 -4207 14459 -4140
rect 12979 -4260 14309 -4207
rect 12979 -5260 13099 -4260
rect 14099 -5260 14309 -4260
rect 12979 -5313 14309 -5260
rect 14397 -5313 14459 -4207
rect 12979 -5380 14459 -5313
rect 14593 -4207 16073 -4140
rect 14593 -4260 15923 -4207
rect 14593 -5260 14713 -4260
rect 15713 -5260 15923 -4260
rect 14593 -5313 15923 -5260
rect 16011 -5313 16073 -4207
rect 14593 -5380 16073 -5313
rect 16207 -4207 17687 -4140
rect 16207 -4260 17537 -4207
rect 16207 -5260 16327 -4260
rect 17327 -5260 17537 -4260
rect 16207 -5313 17537 -5260
rect 17625 -5313 17687 -4207
rect 16207 -5380 17687 -5313
rect -17687 -5567 -16207 -5500
rect -17687 -5620 -16357 -5567
rect -17687 -6620 -17567 -5620
rect -16567 -6620 -16357 -5620
rect -17687 -6673 -16357 -6620
rect -16269 -6673 -16207 -5567
rect -17687 -6740 -16207 -6673
rect -16073 -5567 -14593 -5500
rect -16073 -5620 -14743 -5567
rect -16073 -6620 -15953 -5620
rect -14953 -6620 -14743 -5620
rect -16073 -6673 -14743 -6620
rect -14655 -6673 -14593 -5567
rect -16073 -6740 -14593 -6673
rect -14459 -5567 -12979 -5500
rect -14459 -5620 -13129 -5567
rect -14459 -6620 -14339 -5620
rect -13339 -6620 -13129 -5620
rect -14459 -6673 -13129 -6620
rect -13041 -6673 -12979 -5567
rect -14459 -6740 -12979 -6673
rect -12845 -5567 -11365 -5500
rect -12845 -5620 -11515 -5567
rect -12845 -6620 -12725 -5620
rect -11725 -6620 -11515 -5620
rect -12845 -6673 -11515 -6620
rect -11427 -6673 -11365 -5567
rect -12845 -6740 -11365 -6673
rect -11231 -5567 -9751 -5500
rect -11231 -5620 -9901 -5567
rect -11231 -6620 -11111 -5620
rect -10111 -6620 -9901 -5620
rect -11231 -6673 -9901 -6620
rect -9813 -6673 -9751 -5567
rect -11231 -6740 -9751 -6673
rect -9617 -5567 -8137 -5500
rect -9617 -5620 -8287 -5567
rect -9617 -6620 -9497 -5620
rect -8497 -6620 -8287 -5620
rect -9617 -6673 -8287 -6620
rect -8199 -6673 -8137 -5567
rect -9617 -6740 -8137 -6673
rect -8003 -5567 -6523 -5500
rect -8003 -5620 -6673 -5567
rect -8003 -6620 -7883 -5620
rect -6883 -6620 -6673 -5620
rect -8003 -6673 -6673 -6620
rect -6585 -6673 -6523 -5567
rect -8003 -6740 -6523 -6673
rect -6389 -5567 -4909 -5500
rect -6389 -5620 -5059 -5567
rect -6389 -6620 -6269 -5620
rect -5269 -6620 -5059 -5620
rect -6389 -6673 -5059 -6620
rect -4971 -6673 -4909 -5567
rect -6389 -6740 -4909 -6673
rect -4775 -5567 -3295 -5500
rect -4775 -5620 -3445 -5567
rect -4775 -6620 -4655 -5620
rect -3655 -6620 -3445 -5620
rect -4775 -6673 -3445 -6620
rect -3357 -6673 -3295 -5567
rect -4775 -6740 -3295 -6673
rect -3161 -5567 -1681 -5500
rect -3161 -5620 -1831 -5567
rect -3161 -6620 -3041 -5620
rect -2041 -6620 -1831 -5620
rect -3161 -6673 -1831 -6620
rect -1743 -6673 -1681 -5567
rect -3161 -6740 -1681 -6673
rect -1547 -5567 -67 -5500
rect -1547 -5620 -217 -5567
rect -1547 -6620 -1427 -5620
rect -427 -6620 -217 -5620
rect -1547 -6673 -217 -6620
rect -129 -6673 -67 -5567
rect -1547 -6740 -67 -6673
rect 67 -5567 1547 -5500
rect 67 -5620 1397 -5567
rect 67 -6620 187 -5620
rect 1187 -6620 1397 -5620
rect 67 -6673 1397 -6620
rect 1485 -6673 1547 -5567
rect 67 -6740 1547 -6673
rect 1681 -5567 3161 -5500
rect 1681 -5620 3011 -5567
rect 1681 -6620 1801 -5620
rect 2801 -6620 3011 -5620
rect 1681 -6673 3011 -6620
rect 3099 -6673 3161 -5567
rect 1681 -6740 3161 -6673
rect 3295 -5567 4775 -5500
rect 3295 -5620 4625 -5567
rect 3295 -6620 3415 -5620
rect 4415 -6620 4625 -5620
rect 3295 -6673 4625 -6620
rect 4713 -6673 4775 -5567
rect 3295 -6740 4775 -6673
rect 4909 -5567 6389 -5500
rect 4909 -5620 6239 -5567
rect 4909 -6620 5029 -5620
rect 6029 -6620 6239 -5620
rect 4909 -6673 6239 -6620
rect 6327 -6673 6389 -5567
rect 4909 -6740 6389 -6673
rect 6523 -5567 8003 -5500
rect 6523 -5620 7853 -5567
rect 6523 -6620 6643 -5620
rect 7643 -6620 7853 -5620
rect 6523 -6673 7853 -6620
rect 7941 -6673 8003 -5567
rect 6523 -6740 8003 -6673
rect 8137 -5567 9617 -5500
rect 8137 -5620 9467 -5567
rect 8137 -6620 8257 -5620
rect 9257 -6620 9467 -5620
rect 8137 -6673 9467 -6620
rect 9555 -6673 9617 -5567
rect 8137 -6740 9617 -6673
rect 9751 -5567 11231 -5500
rect 9751 -5620 11081 -5567
rect 9751 -6620 9871 -5620
rect 10871 -6620 11081 -5620
rect 9751 -6673 11081 -6620
rect 11169 -6673 11231 -5567
rect 9751 -6740 11231 -6673
rect 11365 -5567 12845 -5500
rect 11365 -5620 12695 -5567
rect 11365 -6620 11485 -5620
rect 12485 -6620 12695 -5620
rect 11365 -6673 12695 -6620
rect 12783 -6673 12845 -5567
rect 11365 -6740 12845 -6673
rect 12979 -5567 14459 -5500
rect 12979 -5620 14309 -5567
rect 12979 -6620 13099 -5620
rect 14099 -6620 14309 -5620
rect 12979 -6673 14309 -6620
rect 14397 -6673 14459 -5567
rect 12979 -6740 14459 -6673
rect 14593 -5567 16073 -5500
rect 14593 -5620 15923 -5567
rect 14593 -6620 14713 -5620
rect 15713 -6620 15923 -5620
rect 14593 -6673 15923 -6620
rect 16011 -6673 16073 -5567
rect 14593 -6740 16073 -6673
rect 16207 -5567 17687 -5500
rect 16207 -5620 17537 -5567
rect 16207 -6620 16327 -5620
rect 17327 -6620 17537 -5620
rect 16207 -6673 17537 -6620
rect 17625 -6673 17687 -5567
rect 16207 -6740 17687 -6673
rect -17687 -6927 -16207 -6860
rect -17687 -6980 -16357 -6927
rect -17687 -7980 -17567 -6980
rect -16567 -7980 -16357 -6980
rect -17687 -8033 -16357 -7980
rect -16269 -8033 -16207 -6927
rect -17687 -8100 -16207 -8033
rect -16073 -6927 -14593 -6860
rect -16073 -6980 -14743 -6927
rect -16073 -7980 -15953 -6980
rect -14953 -7980 -14743 -6980
rect -16073 -8033 -14743 -7980
rect -14655 -8033 -14593 -6927
rect -16073 -8100 -14593 -8033
rect -14459 -6927 -12979 -6860
rect -14459 -6980 -13129 -6927
rect -14459 -7980 -14339 -6980
rect -13339 -7980 -13129 -6980
rect -14459 -8033 -13129 -7980
rect -13041 -8033 -12979 -6927
rect -14459 -8100 -12979 -8033
rect -12845 -6927 -11365 -6860
rect -12845 -6980 -11515 -6927
rect -12845 -7980 -12725 -6980
rect -11725 -7980 -11515 -6980
rect -12845 -8033 -11515 -7980
rect -11427 -8033 -11365 -6927
rect -12845 -8100 -11365 -8033
rect -11231 -6927 -9751 -6860
rect -11231 -6980 -9901 -6927
rect -11231 -7980 -11111 -6980
rect -10111 -7980 -9901 -6980
rect -11231 -8033 -9901 -7980
rect -9813 -8033 -9751 -6927
rect -11231 -8100 -9751 -8033
rect -9617 -6927 -8137 -6860
rect -9617 -6980 -8287 -6927
rect -9617 -7980 -9497 -6980
rect -8497 -7980 -8287 -6980
rect -9617 -8033 -8287 -7980
rect -8199 -8033 -8137 -6927
rect -9617 -8100 -8137 -8033
rect -8003 -6927 -6523 -6860
rect -8003 -6980 -6673 -6927
rect -8003 -7980 -7883 -6980
rect -6883 -7980 -6673 -6980
rect -8003 -8033 -6673 -7980
rect -6585 -8033 -6523 -6927
rect -8003 -8100 -6523 -8033
rect -6389 -6927 -4909 -6860
rect -6389 -6980 -5059 -6927
rect -6389 -7980 -6269 -6980
rect -5269 -7980 -5059 -6980
rect -6389 -8033 -5059 -7980
rect -4971 -8033 -4909 -6927
rect -6389 -8100 -4909 -8033
rect -4775 -6927 -3295 -6860
rect -4775 -6980 -3445 -6927
rect -4775 -7980 -4655 -6980
rect -3655 -7980 -3445 -6980
rect -4775 -8033 -3445 -7980
rect -3357 -8033 -3295 -6927
rect -4775 -8100 -3295 -8033
rect -3161 -6927 -1681 -6860
rect -3161 -6980 -1831 -6927
rect -3161 -7980 -3041 -6980
rect -2041 -7980 -1831 -6980
rect -3161 -8033 -1831 -7980
rect -1743 -8033 -1681 -6927
rect -3161 -8100 -1681 -8033
rect -1547 -6927 -67 -6860
rect -1547 -6980 -217 -6927
rect -1547 -7980 -1427 -6980
rect -427 -7980 -217 -6980
rect -1547 -8033 -217 -7980
rect -129 -8033 -67 -6927
rect -1547 -8100 -67 -8033
rect 67 -6927 1547 -6860
rect 67 -6980 1397 -6927
rect 67 -7980 187 -6980
rect 1187 -7980 1397 -6980
rect 67 -8033 1397 -7980
rect 1485 -8033 1547 -6927
rect 67 -8100 1547 -8033
rect 1681 -6927 3161 -6860
rect 1681 -6980 3011 -6927
rect 1681 -7980 1801 -6980
rect 2801 -7980 3011 -6980
rect 1681 -8033 3011 -7980
rect 3099 -8033 3161 -6927
rect 1681 -8100 3161 -8033
rect 3295 -6927 4775 -6860
rect 3295 -6980 4625 -6927
rect 3295 -7980 3415 -6980
rect 4415 -7980 4625 -6980
rect 3295 -8033 4625 -7980
rect 4713 -8033 4775 -6927
rect 3295 -8100 4775 -8033
rect 4909 -6927 6389 -6860
rect 4909 -6980 6239 -6927
rect 4909 -7980 5029 -6980
rect 6029 -7980 6239 -6980
rect 4909 -8033 6239 -7980
rect 6327 -8033 6389 -6927
rect 4909 -8100 6389 -8033
rect 6523 -6927 8003 -6860
rect 6523 -6980 7853 -6927
rect 6523 -7980 6643 -6980
rect 7643 -7980 7853 -6980
rect 6523 -8033 7853 -7980
rect 7941 -8033 8003 -6927
rect 6523 -8100 8003 -8033
rect 8137 -6927 9617 -6860
rect 8137 -6980 9467 -6927
rect 8137 -7980 8257 -6980
rect 9257 -7980 9467 -6980
rect 8137 -8033 9467 -7980
rect 9555 -8033 9617 -6927
rect 8137 -8100 9617 -8033
rect 9751 -6927 11231 -6860
rect 9751 -6980 11081 -6927
rect 9751 -7980 9871 -6980
rect 10871 -7980 11081 -6980
rect 9751 -8033 11081 -7980
rect 11169 -8033 11231 -6927
rect 9751 -8100 11231 -8033
rect 11365 -6927 12845 -6860
rect 11365 -6980 12695 -6927
rect 11365 -7980 11485 -6980
rect 12485 -7980 12695 -6980
rect 11365 -8033 12695 -7980
rect 12783 -8033 12845 -6927
rect 11365 -8100 12845 -8033
rect 12979 -6927 14459 -6860
rect 12979 -6980 14309 -6927
rect 12979 -7980 13099 -6980
rect 14099 -7980 14309 -6980
rect 12979 -8033 14309 -7980
rect 14397 -8033 14459 -6927
rect 12979 -8100 14459 -8033
rect 14593 -6927 16073 -6860
rect 14593 -6980 15923 -6927
rect 14593 -7980 14713 -6980
rect 15713 -7980 15923 -6980
rect 14593 -8033 15923 -7980
rect 16011 -8033 16073 -6927
rect 14593 -8100 16073 -8033
rect 16207 -6927 17687 -6860
rect 16207 -6980 17537 -6927
rect 16207 -7980 16327 -6980
rect 17327 -7980 17537 -6980
rect 16207 -8033 17537 -7980
rect 17625 -8033 17687 -6927
rect 16207 -8100 17687 -8033
<< via4 >>
rect -16357 6927 -16269 8033
rect -14743 6927 -14655 8033
rect -13129 6927 -13041 8033
rect -11515 6927 -11427 8033
rect -9901 6927 -9813 8033
rect -8287 6927 -8199 8033
rect -6673 6927 -6585 8033
rect -5059 6927 -4971 8033
rect -3445 6927 -3357 8033
rect -1831 6927 -1743 8033
rect -217 6927 -129 8033
rect 1397 6927 1485 8033
rect 3011 6927 3099 8033
rect 4625 6927 4713 8033
rect 6239 6927 6327 8033
rect 7853 6927 7941 8033
rect 9467 6927 9555 8033
rect 11081 6927 11169 8033
rect 12695 6927 12783 8033
rect 14309 6927 14397 8033
rect 15923 6927 16011 8033
rect 17537 6927 17625 8033
rect -16357 5567 -16269 6673
rect -14743 5567 -14655 6673
rect -13129 5567 -13041 6673
rect -11515 5567 -11427 6673
rect -9901 5567 -9813 6673
rect -8287 5567 -8199 6673
rect -6673 5567 -6585 6673
rect -5059 5567 -4971 6673
rect -3445 5567 -3357 6673
rect -1831 5567 -1743 6673
rect -217 5567 -129 6673
rect 1397 5567 1485 6673
rect 3011 5567 3099 6673
rect 4625 5567 4713 6673
rect 6239 5567 6327 6673
rect 7853 5567 7941 6673
rect 9467 5567 9555 6673
rect 11081 5567 11169 6673
rect 12695 5567 12783 6673
rect 14309 5567 14397 6673
rect 15923 5567 16011 6673
rect 17537 5567 17625 6673
rect -16357 4207 -16269 5313
rect -14743 4207 -14655 5313
rect -13129 4207 -13041 5313
rect -11515 4207 -11427 5313
rect -9901 4207 -9813 5313
rect -8287 4207 -8199 5313
rect -6673 4207 -6585 5313
rect -5059 4207 -4971 5313
rect -3445 4207 -3357 5313
rect -1831 4207 -1743 5313
rect -217 4207 -129 5313
rect 1397 4207 1485 5313
rect 3011 4207 3099 5313
rect 4625 4207 4713 5313
rect 6239 4207 6327 5313
rect 7853 4207 7941 5313
rect 9467 4207 9555 5313
rect 11081 4207 11169 5313
rect 12695 4207 12783 5313
rect 14309 4207 14397 5313
rect 15923 4207 16011 5313
rect 17537 4207 17625 5313
rect -16357 2847 -16269 3953
rect -14743 2847 -14655 3953
rect -13129 2847 -13041 3953
rect -11515 2847 -11427 3953
rect -9901 2847 -9813 3953
rect -8287 2847 -8199 3953
rect -6673 2847 -6585 3953
rect -5059 2847 -4971 3953
rect -3445 2847 -3357 3953
rect -1831 2847 -1743 3953
rect -217 2847 -129 3953
rect 1397 2847 1485 3953
rect 3011 2847 3099 3953
rect 4625 2847 4713 3953
rect 6239 2847 6327 3953
rect 7853 2847 7941 3953
rect 9467 2847 9555 3953
rect 11081 2847 11169 3953
rect 12695 2847 12783 3953
rect 14309 2847 14397 3953
rect 15923 2847 16011 3953
rect 17537 2847 17625 3953
rect -16357 1487 -16269 2593
rect -14743 1487 -14655 2593
rect -13129 1487 -13041 2593
rect -11515 1487 -11427 2593
rect -9901 1487 -9813 2593
rect -8287 1487 -8199 2593
rect -6673 1487 -6585 2593
rect -5059 1487 -4971 2593
rect -3445 1487 -3357 2593
rect -1831 1487 -1743 2593
rect -217 1487 -129 2593
rect 1397 1487 1485 2593
rect 3011 1487 3099 2593
rect 4625 1487 4713 2593
rect 6239 1487 6327 2593
rect 7853 1487 7941 2593
rect 9467 1487 9555 2593
rect 11081 1487 11169 2593
rect 12695 1487 12783 2593
rect 14309 1487 14397 2593
rect 15923 1487 16011 2593
rect 17537 1487 17625 2593
rect -16357 127 -16269 1233
rect -14743 127 -14655 1233
rect -13129 127 -13041 1233
rect -11515 127 -11427 1233
rect -9901 127 -9813 1233
rect -8287 127 -8199 1233
rect -6673 127 -6585 1233
rect -5059 127 -4971 1233
rect -3445 127 -3357 1233
rect -1831 127 -1743 1233
rect -217 127 -129 1233
rect 1397 127 1485 1233
rect 3011 127 3099 1233
rect 4625 127 4713 1233
rect 6239 127 6327 1233
rect 7853 127 7941 1233
rect 9467 127 9555 1233
rect 11081 127 11169 1233
rect 12695 127 12783 1233
rect 14309 127 14397 1233
rect 15923 127 16011 1233
rect 17537 127 17625 1233
rect -16357 -1233 -16269 -127
rect -14743 -1233 -14655 -127
rect -13129 -1233 -13041 -127
rect -11515 -1233 -11427 -127
rect -9901 -1233 -9813 -127
rect -8287 -1233 -8199 -127
rect -6673 -1233 -6585 -127
rect -5059 -1233 -4971 -127
rect -3445 -1233 -3357 -127
rect -1831 -1233 -1743 -127
rect -217 -1233 -129 -127
rect 1397 -1233 1485 -127
rect 3011 -1233 3099 -127
rect 4625 -1233 4713 -127
rect 6239 -1233 6327 -127
rect 7853 -1233 7941 -127
rect 9467 -1233 9555 -127
rect 11081 -1233 11169 -127
rect 12695 -1233 12783 -127
rect 14309 -1233 14397 -127
rect 15923 -1233 16011 -127
rect 17537 -1233 17625 -127
rect -16357 -2593 -16269 -1487
rect -14743 -2593 -14655 -1487
rect -13129 -2593 -13041 -1487
rect -11515 -2593 -11427 -1487
rect -9901 -2593 -9813 -1487
rect -8287 -2593 -8199 -1487
rect -6673 -2593 -6585 -1487
rect -5059 -2593 -4971 -1487
rect -3445 -2593 -3357 -1487
rect -1831 -2593 -1743 -1487
rect -217 -2593 -129 -1487
rect 1397 -2593 1485 -1487
rect 3011 -2593 3099 -1487
rect 4625 -2593 4713 -1487
rect 6239 -2593 6327 -1487
rect 7853 -2593 7941 -1487
rect 9467 -2593 9555 -1487
rect 11081 -2593 11169 -1487
rect 12695 -2593 12783 -1487
rect 14309 -2593 14397 -1487
rect 15923 -2593 16011 -1487
rect 17537 -2593 17625 -1487
rect -16357 -3953 -16269 -2847
rect -14743 -3953 -14655 -2847
rect -13129 -3953 -13041 -2847
rect -11515 -3953 -11427 -2847
rect -9901 -3953 -9813 -2847
rect -8287 -3953 -8199 -2847
rect -6673 -3953 -6585 -2847
rect -5059 -3953 -4971 -2847
rect -3445 -3953 -3357 -2847
rect -1831 -3953 -1743 -2847
rect -217 -3953 -129 -2847
rect 1397 -3953 1485 -2847
rect 3011 -3953 3099 -2847
rect 4625 -3953 4713 -2847
rect 6239 -3953 6327 -2847
rect 7853 -3953 7941 -2847
rect 9467 -3953 9555 -2847
rect 11081 -3953 11169 -2847
rect 12695 -3953 12783 -2847
rect 14309 -3953 14397 -2847
rect 15923 -3953 16011 -2847
rect 17537 -3953 17625 -2847
rect -16357 -5313 -16269 -4207
rect -14743 -5313 -14655 -4207
rect -13129 -5313 -13041 -4207
rect -11515 -5313 -11427 -4207
rect -9901 -5313 -9813 -4207
rect -8287 -5313 -8199 -4207
rect -6673 -5313 -6585 -4207
rect -5059 -5313 -4971 -4207
rect -3445 -5313 -3357 -4207
rect -1831 -5313 -1743 -4207
rect -217 -5313 -129 -4207
rect 1397 -5313 1485 -4207
rect 3011 -5313 3099 -4207
rect 4625 -5313 4713 -4207
rect 6239 -5313 6327 -4207
rect 7853 -5313 7941 -4207
rect 9467 -5313 9555 -4207
rect 11081 -5313 11169 -4207
rect 12695 -5313 12783 -4207
rect 14309 -5313 14397 -4207
rect 15923 -5313 16011 -4207
rect 17537 -5313 17625 -4207
rect -16357 -6673 -16269 -5567
rect -14743 -6673 -14655 -5567
rect -13129 -6673 -13041 -5567
rect -11515 -6673 -11427 -5567
rect -9901 -6673 -9813 -5567
rect -8287 -6673 -8199 -5567
rect -6673 -6673 -6585 -5567
rect -5059 -6673 -4971 -5567
rect -3445 -6673 -3357 -5567
rect -1831 -6673 -1743 -5567
rect -217 -6673 -129 -5567
rect 1397 -6673 1485 -5567
rect 3011 -6673 3099 -5567
rect 4625 -6673 4713 -5567
rect 6239 -6673 6327 -5567
rect 7853 -6673 7941 -5567
rect 9467 -6673 9555 -5567
rect 11081 -6673 11169 -5567
rect 12695 -6673 12783 -5567
rect 14309 -6673 14397 -5567
rect 15923 -6673 16011 -5567
rect 17537 -6673 17625 -5567
rect -16357 -8033 -16269 -6927
rect -14743 -8033 -14655 -6927
rect -13129 -8033 -13041 -6927
rect -11515 -8033 -11427 -6927
rect -9901 -8033 -9813 -6927
rect -8287 -8033 -8199 -6927
rect -6673 -8033 -6585 -6927
rect -5059 -8033 -4971 -6927
rect -3445 -8033 -3357 -6927
rect -1831 -8033 -1743 -6927
rect -217 -8033 -129 -6927
rect 1397 -8033 1485 -6927
rect 3011 -8033 3099 -6927
rect 4625 -8033 4713 -6927
rect 6239 -8033 6327 -6927
rect 7853 -8033 7941 -6927
rect 9467 -8033 9555 -6927
rect 11081 -8033 11169 -6927
rect 12695 -8033 12783 -6927
rect 14309 -8033 14397 -6927
rect 15923 -8033 16011 -6927
rect 17537 -8033 17625 -6927
<< metal5 >>
rect -17173 7900 -16961 8160
rect -16419 8033 -16207 8160
rect -17173 6540 -16961 7060
rect -16419 6927 -16357 8033
rect -16269 6927 -16207 8033
rect -15559 7900 -15347 8160
rect -14805 8033 -14593 8160
rect -16419 6673 -16207 6927
rect -17173 5180 -16961 5700
rect -16419 5567 -16357 6673
rect -16269 5567 -16207 6673
rect -15559 6540 -15347 7060
rect -14805 6927 -14743 8033
rect -14655 6927 -14593 8033
rect -13945 7900 -13733 8160
rect -13191 8033 -12979 8160
rect -14805 6673 -14593 6927
rect -16419 5313 -16207 5567
rect -17173 3820 -16961 4340
rect -16419 4207 -16357 5313
rect -16269 4207 -16207 5313
rect -15559 5180 -15347 5700
rect -14805 5567 -14743 6673
rect -14655 5567 -14593 6673
rect -13945 6540 -13733 7060
rect -13191 6927 -13129 8033
rect -13041 6927 -12979 8033
rect -12331 7900 -12119 8160
rect -11577 8033 -11365 8160
rect -13191 6673 -12979 6927
rect -14805 5313 -14593 5567
rect -16419 3953 -16207 4207
rect -17173 2460 -16961 2980
rect -16419 2847 -16357 3953
rect -16269 2847 -16207 3953
rect -15559 3820 -15347 4340
rect -14805 4207 -14743 5313
rect -14655 4207 -14593 5313
rect -13945 5180 -13733 5700
rect -13191 5567 -13129 6673
rect -13041 5567 -12979 6673
rect -12331 6540 -12119 7060
rect -11577 6927 -11515 8033
rect -11427 6927 -11365 8033
rect -10717 7900 -10505 8160
rect -9963 8033 -9751 8160
rect -11577 6673 -11365 6927
rect -13191 5313 -12979 5567
rect -14805 3953 -14593 4207
rect -16419 2593 -16207 2847
rect -17173 1100 -16961 1620
rect -16419 1487 -16357 2593
rect -16269 1487 -16207 2593
rect -15559 2460 -15347 2980
rect -14805 2847 -14743 3953
rect -14655 2847 -14593 3953
rect -13945 3820 -13733 4340
rect -13191 4207 -13129 5313
rect -13041 4207 -12979 5313
rect -12331 5180 -12119 5700
rect -11577 5567 -11515 6673
rect -11427 5567 -11365 6673
rect -10717 6540 -10505 7060
rect -9963 6927 -9901 8033
rect -9813 6927 -9751 8033
rect -9103 7900 -8891 8160
rect -8349 8033 -8137 8160
rect -9963 6673 -9751 6927
rect -11577 5313 -11365 5567
rect -13191 3953 -12979 4207
rect -14805 2593 -14593 2847
rect -16419 1233 -16207 1487
rect -17173 -260 -16961 260
rect -16419 127 -16357 1233
rect -16269 127 -16207 1233
rect -15559 1100 -15347 1620
rect -14805 1487 -14743 2593
rect -14655 1487 -14593 2593
rect -13945 2460 -13733 2980
rect -13191 2847 -13129 3953
rect -13041 2847 -12979 3953
rect -12331 3820 -12119 4340
rect -11577 4207 -11515 5313
rect -11427 4207 -11365 5313
rect -10717 5180 -10505 5700
rect -9963 5567 -9901 6673
rect -9813 5567 -9751 6673
rect -9103 6540 -8891 7060
rect -8349 6927 -8287 8033
rect -8199 6927 -8137 8033
rect -7489 7900 -7277 8160
rect -6735 8033 -6523 8160
rect -8349 6673 -8137 6927
rect -9963 5313 -9751 5567
rect -11577 3953 -11365 4207
rect -13191 2593 -12979 2847
rect -14805 1233 -14593 1487
rect -16419 -127 -16207 127
rect -17173 -1620 -16961 -1100
rect -16419 -1233 -16357 -127
rect -16269 -1233 -16207 -127
rect -15559 -260 -15347 260
rect -14805 127 -14743 1233
rect -14655 127 -14593 1233
rect -13945 1100 -13733 1620
rect -13191 1487 -13129 2593
rect -13041 1487 -12979 2593
rect -12331 2460 -12119 2980
rect -11577 2847 -11515 3953
rect -11427 2847 -11365 3953
rect -10717 3820 -10505 4340
rect -9963 4207 -9901 5313
rect -9813 4207 -9751 5313
rect -9103 5180 -8891 5700
rect -8349 5567 -8287 6673
rect -8199 5567 -8137 6673
rect -7489 6540 -7277 7060
rect -6735 6927 -6673 8033
rect -6585 6927 -6523 8033
rect -5875 7900 -5663 8160
rect -5121 8033 -4909 8160
rect -6735 6673 -6523 6927
rect -8349 5313 -8137 5567
rect -9963 3953 -9751 4207
rect -11577 2593 -11365 2847
rect -13191 1233 -12979 1487
rect -14805 -127 -14593 127
rect -16419 -1487 -16207 -1233
rect -17173 -2980 -16961 -2460
rect -16419 -2593 -16357 -1487
rect -16269 -2593 -16207 -1487
rect -15559 -1620 -15347 -1100
rect -14805 -1233 -14743 -127
rect -14655 -1233 -14593 -127
rect -13945 -260 -13733 260
rect -13191 127 -13129 1233
rect -13041 127 -12979 1233
rect -12331 1100 -12119 1620
rect -11577 1487 -11515 2593
rect -11427 1487 -11365 2593
rect -10717 2460 -10505 2980
rect -9963 2847 -9901 3953
rect -9813 2847 -9751 3953
rect -9103 3820 -8891 4340
rect -8349 4207 -8287 5313
rect -8199 4207 -8137 5313
rect -7489 5180 -7277 5700
rect -6735 5567 -6673 6673
rect -6585 5567 -6523 6673
rect -5875 6540 -5663 7060
rect -5121 6927 -5059 8033
rect -4971 6927 -4909 8033
rect -4261 7900 -4049 8160
rect -3507 8033 -3295 8160
rect -5121 6673 -4909 6927
rect -6735 5313 -6523 5567
rect -8349 3953 -8137 4207
rect -9963 2593 -9751 2847
rect -11577 1233 -11365 1487
rect -13191 -127 -12979 127
rect -14805 -1487 -14593 -1233
rect -16419 -2847 -16207 -2593
rect -17173 -4340 -16961 -3820
rect -16419 -3953 -16357 -2847
rect -16269 -3953 -16207 -2847
rect -15559 -2980 -15347 -2460
rect -14805 -2593 -14743 -1487
rect -14655 -2593 -14593 -1487
rect -13945 -1620 -13733 -1100
rect -13191 -1233 -13129 -127
rect -13041 -1233 -12979 -127
rect -12331 -260 -12119 260
rect -11577 127 -11515 1233
rect -11427 127 -11365 1233
rect -10717 1100 -10505 1620
rect -9963 1487 -9901 2593
rect -9813 1487 -9751 2593
rect -9103 2460 -8891 2980
rect -8349 2847 -8287 3953
rect -8199 2847 -8137 3953
rect -7489 3820 -7277 4340
rect -6735 4207 -6673 5313
rect -6585 4207 -6523 5313
rect -5875 5180 -5663 5700
rect -5121 5567 -5059 6673
rect -4971 5567 -4909 6673
rect -4261 6540 -4049 7060
rect -3507 6927 -3445 8033
rect -3357 6927 -3295 8033
rect -2647 7900 -2435 8160
rect -1893 8033 -1681 8160
rect -3507 6673 -3295 6927
rect -5121 5313 -4909 5567
rect -6735 3953 -6523 4207
rect -8349 2593 -8137 2847
rect -9963 1233 -9751 1487
rect -11577 -127 -11365 127
rect -13191 -1487 -12979 -1233
rect -14805 -2847 -14593 -2593
rect -16419 -4207 -16207 -3953
rect -17173 -5700 -16961 -5180
rect -16419 -5313 -16357 -4207
rect -16269 -5313 -16207 -4207
rect -15559 -4340 -15347 -3820
rect -14805 -3953 -14743 -2847
rect -14655 -3953 -14593 -2847
rect -13945 -2980 -13733 -2460
rect -13191 -2593 -13129 -1487
rect -13041 -2593 -12979 -1487
rect -12331 -1620 -12119 -1100
rect -11577 -1233 -11515 -127
rect -11427 -1233 -11365 -127
rect -10717 -260 -10505 260
rect -9963 127 -9901 1233
rect -9813 127 -9751 1233
rect -9103 1100 -8891 1620
rect -8349 1487 -8287 2593
rect -8199 1487 -8137 2593
rect -7489 2460 -7277 2980
rect -6735 2847 -6673 3953
rect -6585 2847 -6523 3953
rect -5875 3820 -5663 4340
rect -5121 4207 -5059 5313
rect -4971 4207 -4909 5313
rect -4261 5180 -4049 5700
rect -3507 5567 -3445 6673
rect -3357 5567 -3295 6673
rect -2647 6540 -2435 7060
rect -1893 6927 -1831 8033
rect -1743 6927 -1681 8033
rect -1033 7900 -821 8160
rect -279 8033 -67 8160
rect -1893 6673 -1681 6927
rect -3507 5313 -3295 5567
rect -5121 3953 -4909 4207
rect -6735 2593 -6523 2847
rect -8349 1233 -8137 1487
rect -9963 -127 -9751 127
rect -11577 -1487 -11365 -1233
rect -13191 -2847 -12979 -2593
rect -14805 -4207 -14593 -3953
rect -16419 -5567 -16207 -5313
rect -17173 -7060 -16961 -6540
rect -16419 -6673 -16357 -5567
rect -16269 -6673 -16207 -5567
rect -15559 -5700 -15347 -5180
rect -14805 -5313 -14743 -4207
rect -14655 -5313 -14593 -4207
rect -13945 -4340 -13733 -3820
rect -13191 -3953 -13129 -2847
rect -13041 -3953 -12979 -2847
rect -12331 -2980 -12119 -2460
rect -11577 -2593 -11515 -1487
rect -11427 -2593 -11365 -1487
rect -10717 -1620 -10505 -1100
rect -9963 -1233 -9901 -127
rect -9813 -1233 -9751 -127
rect -9103 -260 -8891 260
rect -8349 127 -8287 1233
rect -8199 127 -8137 1233
rect -7489 1100 -7277 1620
rect -6735 1487 -6673 2593
rect -6585 1487 -6523 2593
rect -5875 2460 -5663 2980
rect -5121 2847 -5059 3953
rect -4971 2847 -4909 3953
rect -4261 3820 -4049 4340
rect -3507 4207 -3445 5313
rect -3357 4207 -3295 5313
rect -2647 5180 -2435 5700
rect -1893 5567 -1831 6673
rect -1743 5567 -1681 6673
rect -1033 6540 -821 7060
rect -279 6927 -217 8033
rect -129 6927 -67 8033
rect 581 7900 793 8160
rect 1335 8033 1547 8160
rect -279 6673 -67 6927
rect -1893 5313 -1681 5567
rect -3507 3953 -3295 4207
rect -5121 2593 -4909 2847
rect -6735 1233 -6523 1487
rect -8349 -127 -8137 127
rect -9963 -1487 -9751 -1233
rect -11577 -2847 -11365 -2593
rect -13191 -4207 -12979 -3953
rect -14805 -5567 -14593 -5313
rect -16419 -6927 -16207 -6673
rect -17173 -8160 -16961 -7900
rect -16419 -8033 -16357 -6927
rect -16269 -8033 -16207 -6927
rect -15559 -7060 -15347 -6540
rect -14805 -6673 -14743 -5567
rect -14655 -6673 -14593 -5567
rect -13945 -5700 -13733 -5180
rect -13191 -5313 -13129 -4207
rect -13041 -5313 -12979 -4207
rect -12331 -4340 -12119 -3820
rect -11577 -3953 -11515 -2847
rect -11427 -3953 -11365 -2847
rect -10717 -2980 -10505 -2460
rect -9963 -2593 -9901 -1487
rect -9813 -2593 -9751 -1487
rect -9103 -1620 -8891 -1100
rect -8349 -1233 -8287 -127
rect -8199 -1233 -8137 -127
rect -7489 -260 -7277 260
rect -6735 127 -6673 1233
rect -6585 127 -6523 1233
rect -5875 1100 -5663 1620
rect -5121 1487 -5059 2593
rect -4971 1487 -4909 2593
rect -4261 2460 -4049 2980
rect -3507 2847 -3445 3953
rect -3357 2847 -3295 3953
rect -2647 3820 -2435 4340
rect -1893 4207 -1831 5313
rect -1743 4207 -1681 5313
rect -1033 5180 -821 5700
rect -279 5567 -217 6673
rect -129 5567 -67 6673
rect 581 6540 793 7060
rect 1335 6927 1397 8033
rect 1485 6927 1547 8033
rect 2195 7900 2407 8160
rect 2949 8033 3161 8160
rect 1335 6673 1547 6927
rect -279 5313 -67 5567
rect -1893 3953 -1681 4207
rect -3507 2593 -3295 2847
rect -5121 1233 -4909 1487
rect -6735 -127 -6523 127
rect -8349 -1487 -8137 -1233
rect -9963 -2847 -9751 -2593
rect -11577 -4207 -11365 -3953
rect -13191 -5567 -12979 -5313
rect -14805 -6927 -14593 -6673
rect -16419 -8160 -16207 -8033
rect -15559 -8160 -15347 -7900
rect -14805 -8033 -14743 -6927
rect -14655 -8033 -14593 -6927
rect -13945 -7060 -13733 -6540
rect -13191 -6673 -13129 -5567
rect -13041 -6673 -12979 -5567
rect -12331 -5700 -12119 -5180
rect -11577 -5313 -11515 -4207
rect -11427 -5313 -11365 -4207
rect -10717 -4340 -10505 -3820
rect -9963 -3953 -9901 -2847
rect -9813 -3953 -9751 -2847
rect -9103 -2980 -8891 -2460
rect -8349 -2593 -8287 -1487
rect -8199 -2593 -8137 -1487
rect -7489 -1620 -7277 -1100
rect -6735 -1233 -6673 -127
rect -6585 -1233 -6523 -127
rect -5875 -260 -5663 260
rect -5121 127 -5059 1233
rect -4971 127 -4909 1233
rect -4261 1100 -4049 1620
rect -3507 1487 -3445 2593
rect -3357 1487 -3295 2593
rect -2647 2460 -2435 2980
rect -1893 2847 -1831 3953
rect -1743 2847 -1681 3953
rect -1033 3820 -821 4340
rect -279 4207 -217 5313
rect -129 4207 -67 5313
rect 581 5180 793 5700
rect 1335 5567 1397 6673
rect 1485 5567 1547 6673
rect 2195 6540 2407 7060
rect 2949 6927 3011 8033
rect 3099 6927 3161 8033
rect 3809 7900 4021 8160
rect 4563 8033 4775 8160
rect 2949 6673 3161 6927
rect 1335 5313 1547 5567
rect -279 3953 -67 4207
rect -1893 2593 -1681 2847
rect -3507 1233 -3295 1487
rect -5121 -127 -4909 127
rect -6735 -1487 -6523 -1233
rect -8349 -2847 -8137 -2593
rect -9963 -4207 -9751 -3953
rect -11577 -5567 -11365 -5313
rect -13191 -6927 -12979 -6673
rect -14805 -8160 -14593 -8033
rect -13945 -8160 -13733 -7900
rect -13191 -8033 -13129 -6927
rect -13041 -8033 -12979 -6927
rect -12331 -7060 -12119 -6540
rect -11577 -6673 -11515 -5567
rect -11427 -6673 -11365 -5567
rect -10717 -5700 -10505 -5180
rect -9963 -5313 -9901 -4207
rect -9813 -5313 -9751 -4207
rect -9103 -4340 -8891 -3820
rect -8349 -3953 -8287 -2847
rect -8199 -3953 -8137 -2847
rect -7489 -2980 -7277 -2460
rect -6735 -2593 -6673 -1487
rect -6585 -2593 -6523 -1487
rect -5875 -1620 -5663 -1100
rect -5121 -1233 -5059 -127
rect -4971 -1233 -4909 -127
rect -4261 -260 -4049 260
rect -3507 127 -3445 1233
rect -3357 127 -3295 1233
rect -2647 1100 -2435 1620
rect -1893 1487 -1831 2593
rect -1743 1487 -1681 2593
rect -1033 2460 -821 2980
rect -279 2847 -217 3953
rect -129 2847 -67 3953
rect 581 3820 793 4340
rect 1335 4207 1397 5313
rect 1485 4207 1547 5313
rect 2195 5180 2407 5700
rect 2949 5567 3011 6673
rect 3099 5567 3161 6673
rect 3809 6540 4021 7060
rect 4563 6927 4625 8033
rect 4713 6927 4775 8033
rect 5423 7900 5635 8160
rect 6177 8033 6389 8160
rect 4563 6673 4775 6927
rect 2949 5313 3161 5567
rect 1335 3953 1547 4207
rect -279 2593 -67 2847
rect -1893 1233 -1681 1487
rect -3507 -127 -3295 127
rect -5121 -1487 -4909 -1233
rect -6735 -2847 -6523 -2593
rect -8349 -4207 -8137 -3953
rect -9963 -5567 -9751 -5313
rect -11577 -6927 -11365 -6673
rect -13191 -8160 -12979 -8033
rect -12331 -8160 -12119 -7900
rect -11577 -8033 -11515 -6927
rect -11427 -8033 -11365 -6927
rect -10717 -7060 -10505 -6540
rect -9963 -6673 -9901 -5567
rect -9813 -6673 -9751 -5567
rect -9103 -5700 -8891 -5180
rect -8349 -5313 -8287 -4207
rect -8199 -5313 -8137 -4207
rect -7489 -4340 -7277 -3820
rect -6735 -3953 -6673 -2847
rect -6585 -3953 -6523 -2847
rect -5875 -2980 -5663 -2460
rect -5121 -2593 -5059 -1487
rect -4971 -2593 -4909 -1487
rect -4261 -1620 -4049 -1100
rect -3507 -1233 -3445 -127
rect -3357 -1233 -3295 -127
rect -2647 -260 -2435 260
rect -1893 127 -1831 1233
rect -1743 127 -1681 1233
rect -1033 1100 -821 1620
rect -279 1487 -217 2593
rect -129 1487 -67 2593
rect 581 2460 793 2980
rect 1335 2847 1397 3953
rect 1485 2847 1547 3953
rect 2195 3820 2407 4340
rect 2949 4207 3011 5313
rect 3099 4207 3161 5313
rect 3809 5180 4021 5700
rect 4563 5567 4625 6673
rect 4713 5567 4775 6673
rect 5423 6540 5635 7060
rect 6177 6927 6239 8033
rect 6327 6927 6389 8033
rect 7037 7900 7249 8160
rect 7791 8033 8003 8160
rect 6177 6673 6389 6927
rect 4563 5313 4775 5567
rect 2949 3953 3161 4207
rect 1335 2593 1547 2847
rect -279 1233 -67 1487
rect -1893 -127 -1681 127
rect -3507 -1487 -3295 -1233
rect -5121 -2847 -4909 -2593
rect -6735 -4207 -6523 -3953
rect -8349 -5567 -8137 -5313
rect -9963 -6927 -9751 -6673
rect -11577 -8160 -11365 -8033
rect -10717 -8160 -10505 -7900
rect -9963 -8033 -9901 -6927
rect -9813 -8033 -9751 -6927
rect -9103 -7060 -8891 -6540
rect -8349 -6673 -8287 -5567
rect -8199 -6673 -8137 -5567
rect -7489 -5700 -7277 -5180
rect -6735 -5313 -6673 -4207
rect -6585 -5313 -6523 -4207
rect -5875 -4340 -5663 -3820
rect -5121 -3953 -5059 -2847
rect -4971 -3953 -4909 -2847
rect -4261 -2980 -4049 -2460
rect -3507 -2593 -3445 -1487
rect -3357 -2593 -3295 -1487
rect -2647 -1620 -2435 -1100
rect -1893 -1233 -1831 -127
rect -1743 -1233 -1681 -127
rect -1033 -260 -821 260
rect -279 127 -217 1233
rect -129 127 -67 1233
rect 581 1100 793 1620
rect 1335 1487 1397 2593
rect 1485 1487 1547 2593
rect 2195 2460 2407 2980
rect 2949 2847 3011 3953
rect 3099 2847 3161 3953
rect 3809 3820 4021 4340
rect 4563 4207 4625 5313
rect 4713 4207 4775 5313
rect 5423 5180 5635 5700
rect 6177 5567 6239 6673
rect 6327 5567 6389 6673
rect 7037 6540 7249 7060
rect 7791 6927 7853 8033
rect 7941 6927 8003 8033
rect 8651 7900 8863 8160
rect 9405 8033 9617 8160
rect 7791 6673 8003 6927
rect 6177 5313 6389 5567
rect 4563 3953 4775 4207
rect 2949 2593 3161 2847
rect 1335 1233 1547 1487
rect -279 -127 -67 127
rect -1893 -1487 -1681 -1233
rect -3507 -2847 -3295 -2593
rect -5121 -4207 -4909 -3953
rect -6735 -5567 -6523 -5313
rect -8349 -6927 -8137 -6673
rect -9963 -8160 -9751 -8033
rect -9103 -8160 -8891 -7900
rect -8349 -8033 -8287 -6927
rect -8199 -8033 -8137 -6927
rect -7489 -7060 -7277 -6540
rect -6735 -6673 -6673 -5567
rect -6585 -6673 -6523 -5567
rect -5875 -5700 -5663 -5180
rect -5121 -5313 -5059 -4207
rect -4971 -5313 -4909 -4207
rect -4261 -4340 -4049 -3820
rect -3507 -3953 -3445 -2847
rect -3357 -3953 -3295 -2847
rect -2647 -2980 -2435 -2460
rect -1893 -2593 -1831 -1487
rect -1743 -2593 -1681 -1487
rect -1033 -1620 -821 -1100
rect -279 -1233 -217 -127
rect -129 -1233 -67 -127
rect 581 -260 793 260
rect 1335 127 1397 1233
rect 1485 127 1547 1233
rect 2195 1100 2407 1620
rect 2949 1487 3011 2593
rect 3099 1487 3161 2593
rect 3809 2460 4021 2980
rect 4563 2847 4625 3953
rect 4713 2847 4775 3953
rect 5423 3820 5635 4340
rect 6177 4207 6239 5313
rect 6327 4207 6389 5313
rect 7037 5180 7249 5700
rect 7791 5567 7853 6673
rect 7941 5567 8003 6673
rect 8651 6540 8863 7060
rect 9405 6927 9467 8033
rect 9555 6927 9617 8033
rect 10265 7900 10477 8160
rect 11019 8033 11231 8160
rect 9405 6673 9617 6927
rect 7791 5313 8003 5567
rect 6177 3953 6389 4207
rect 4563 2593 4775 2847
rect 2949 1233 3161 1487
rect 1335 -127 1547 127
rect -279 -1487 -67 -1233
rect -1893 -2847 -1681 -2593
rect -3507 -4207 -3295 -3953
rect -5121 -5567 -4909 -5313
rect -6735 -6927 -6523 -6673
rect -8349 -8160 -8137 -8033
rect -7489 -8160 -7277 -7900
rect -6735 -8033 -6673 -6927
rect -6585 -8033 -6523 -6927
rect -5875 -7060 -5663 -6540
rect -5121 -6673 -5059 -5567
rect -4971 -6673 -4909 -5567
rect -4261 -5700 -4049 -5180
rect -3507 -5313 -3445 -4207
rect -3357 -5313 -3295 -4207
rect -2647 -4340 -2435 -3820
rect -1893 -3953 -1831 -2847
rect -1743 -3953 -1681 -2847
rect -1033 -2980 -821 -2460
rect -279 -2593 -217 -1487
rect -129 -2593 -67 -1487
rect 581 -1620 793 -1100
rect 1335 -1233 1397 -127
rect 1485 -1233 1547 -127
rect 2195 -260 2407 260
rect 2949 127 3011 1233
rect 3099 127 3161 1233
rect 3809 1100 4021 1620
rect 4563 1487 4625 2593
rect 4713 1487 4775 2593
rect 5423 2460 5635 2980
rect 6177 2847 6239 3953
rect 6327 2847 6389 3953
rect 7037 3820 7249 4340
rect 7791 4207 7853 5313
rect 7941 4207 8003 5313
rect 8651 5180 8863 5700
rect 9405 5567 9467 6673
rect 9555 5567 9617 6673
rect 10265 6540 10477 7060
rect 11019 6927 11081 8033
rect 11169 6927 11231 8033
rect 11879 7900 12091 8160
rect 12633 8033 12845 8160
rect 11019 6673 11231 6927
rect 9405 5313 9617 5567
rect 7791 3953 8003 4207
rect 6177 2593 6389 2847
rect 4563 1233 4775 1487
rect 2949 -127 3161 127
rect 1335 -1487 1547 -1233
rect -279 -2847 -67 -2593
rect -1893 -4207 -1681 -3953
rect -3507 -5567 -3295 -5313
rect -5121 -6927 -4909 -6673
rect -6735 -8160 -6523 -8033
rect -5875 -8160 -5663 -7900
rect -5121 -8033 -5059 -6927
rect -4971 -8033 -4909 -6927
rect -4261 -7060 -4049 -6540
rect -3507 -6673 -3445 -5567
rect -3357 -6673 -3295 -5567
rect -2647 -5700 -2435 -5180
rect -1893 -5313 -1831 -4207
rect -1743 -5313 -1681 -4207
rect -1033 -4340 -821 -3820
rect -279 -3953 -217 -2847
rect -129 -3953 -67 -2847
rect 581 -2980 793 -2460
rect 1335 -2593 1397 -1487
rect 1485 -2593 1547 -1487
rect 2195 -1620 2407 -1100
rect 2949 -1233 3011 -127
rect 3099 -1233 3161 -127
rect 3809 -260 4021 260
rect 4563 127 4625 1233
rect 4713 127 4775 1233
rect 5423 1100 5635 1620
rect 6177 1487 6239 2593
rect 6327 1487 6389 2593
rect 7037 2460 7249 2980
rect 7791 2847 7853 3953
rect 7941 2847 8003 3953
rect 8651 3820 8863 4340
rect 9405 4207 9467 5313
rect 9555 4207 9617 5313
rect 10265 5180 10477 5700
rect 11019 5567 11081 6673
rect 11169 5567 11231 6673
rect 11879 6540 12091 7060
rect 12633 6927 12695 8033
rect 12783 6927 12845 8033
rect 13493 7900 13705 8160
rect 14247 8033 14459 8160
rect 12633 6673 12845 6927
rect 11019 5313 11231 5567
rect 9405 3953 9617 4207
rect 7791 2593 8003 2847
rect 6177 1233 6389 1487
rect 4563 -127 4775 127
rect 2949 -1487 3161 -1233
rect 1335 -2847 1547 -2593
rect -279 -4207 -67 -3953
rect -1893 -5567 -1681 -5313
rect -3507 -6927 -3295 -6673
rect -5121 -8160 -4909 -8033
rect -4261 -8160 -4049 -7900
rect -3507 -8033 -3445 -6927
rect -3357 -8033 -3295 -6927
rect -2647 -7060 -2435 -6540
rect -1893 -6673 -1831 -5567
rect -1743 -6673 -1681 -5567
rect -1033 -5700 -821 -5180
rect -279 -5313 -217 -4207
rect -129 -5313 -67 -4207
rect 581 -4340 793 -3820
rect 1335 -3953 1397 -2847
rect 1485 -3953 1547 -2847
rect 2195 -2980 2407 -2460
rect 2949 -2593 3011 -1487
rect 3099 -2593 3161 -1487
rect 3809 -1620 4021 -1100
rect 4563 -1233 4625 -127
rect 4713 -1233 4775 -127
rect 5423 -260 5635 260
rect 6177 127 6239 1233
rect 6327 127 6389 1233
rect 7037 1100 7249 1620
rect 7791 1487 7853 2593
rect 7941 1487 8003 2593
rect 8651 2460 8863 2980
rect 9405 2847 9467 3953
rect 9555 2847 9617 3953
rect 10265 3820 10477 4340
rect 11019 4207 11081 5313
rect 11169 4207 11231 5313
rect 11879 5180 12091 5700
rect 12633 5567 12695 6673
rect 12783 5567 12845 6673
rect 13493 6540 13705 7060
rect 14247 6927 14309 8033
rect 14397 6927 14459 8033
rect 15107 7900 15319 8160
rect 15861 8033 16073 8160
rect 14247 6673 14459 6927
rect 12633 5313 12845 5567
rect 11019 3953 11231 4207
rect 9405 2593 9617 2847
rect 7791 1233 8003 1487
rect 6177 -127 6389 127
rect 4563 -1487 4775 -1233
rect 2949 -2847 3161 -2593
rect 1335 -4207 1547 -3953
rect -279 -5567 -67 -5313
rect -1893 -6927 -1681 -6673
rect -3507 -8160 -3295 -8033
rect -2647 -8160 -2435 -7900
rect -1893 -8033 -1831 -6927
rect -1743 -8033 -1681 -6927
rect -1033 -7060 -821 -6540
rect -279 -6673 -217 -5567
rect -129 -6673 -67 -5567
rect 581 -5700 793 -5180
rect 1335 -5313 1397 -4207
rect 1485 -5313 1547 -4207
rect 2195 -4340 2407 -3820
rect 2949 -3953 3011 -2847
rect 3099 -3953 3161 -2847
rect 3809 -2980 4021 -2460
rect 4563 -2593 4625 -1487
rect 4713 -2593 4775 -1487
rect 5423 -1620 5635 -1100
rect 6177 -1233 6239 -127
rect 6327 -1233 6389 -127
rect 7037 -260 7249 260
rect 7791 127 7853 1233
rect 7941 127 8003 1233
rect 8651 1100 8863 1620
rect 9405 1487 9467 2593
rect 9555 1487 9617 2593
rect 10265 2460 10477 2980
rect 11019 2847 11081 3953
rect 11169 2847 11231 3953
rect 11879 3820 12091 4340
rect 12633 4207 12695 5313
rect 12783 4207 12845 5313
rect 13493 5180 13705 5700
rect 14247 5567 14309 6673
rect 14397 5567 14459 6673
rect 15107 6540 15319 7060
rect 15861 6927 15923 8033
rect 16011 6927 16073 8033
rect 16721 7900 16933 8160
rect 17475 8033 17687 8160
rect 15861 6673 16073 6927
rect 14247 5313 14459 5567
rect 12633 3953 12845 4207
rect 11019 2593 11231 2847
rect 9405 1233 9617 1487
rect 7791 -127 8003 127
rect 6177 -1487 6389 -1233
rect 4563 -2847 4775 -2593
rect 2949 -4207 3161 -3953
rect 1335 -5567 1547 -5313
rect -279 -6927 -67 -6673
rect -1893 -8160 -1681 -8033
rect -1033 -8160 -821 -7900
rect -279 -8033 -217 -6927
rect -129 -8033 -67 -6927
rect 581 -7060 793 -6540
rect 1335 -6673 1397 -5567
rect 1485 -6673 1547 -5567
rect 2195 -5700 2407 -5180
rect 2949 -5313 3011 -4207
rect 3099 -5313 3161 -4207
rect 3809 -4340 4021 -3820
rect 4563 -3953 4625 -2847
rect 4713 -3953 4775 -2847
rect 5423 -2980 5635 -2460
rect 6177 -2593 6239 -1487
rect 6327 -2593 6389 -1487
rect 7037 -1620 7249 -1100
rect 7791 -1233 7853 -127
rect 7941 -1233 8003 -127
rect 8651 -260 8863 260
rect 9405 127 9467 1233
rect 9555 127 9617 1233
rect 10265 1100 10477 1620
rect 11019 1487 11081 2593
rect 11169 1487 11231 2593
rect 11879 2460 12091 2980
rect 12633 2847 12695 3953
rect 12783 2847 12845 3953
rect 13493 3820 13705 4340
rect 14247 4207 14309 5313
rect 14397 4207 14459 5313
rect 15107 5180 15319 5700
rect 15861 5567 15923 6673
rect 16011 5567 16073 6673
rect 16721 6540 16933 7060
rect 17475 6927 17537 8033
rect 17625 6927 17687 8033
rect 17475 6673 17687 6927
rect 15861 5313 16073 5567
rect 14247 3953 14459 4207
rect 12633 2593 12845 2847
rect 11019 1233 11231 1487
rect 9405 -127 9617 127
rect 7791 -1487 8003 -1233
rect 6177 -2847 6389 -2593
rect 4563 -4207 4775 -3953
rect 2949 -5567 3161 -5313
rect 1335 -6927 1547 -6673
rect -279 -8160 -67 -8033
rect 581 -8160 793 -7900
rect 1335 -8033 1397 -6927
rect 1485 -8033 1547 -6927
rect 2195 -7060 2407 -6540
rect 2949 -6673 3011 -5567
rect 3099 -6673 3161 -5567
rect 3809 -5700 4021 -5180
rect 4563 -5313 4625 -4207
rect 4713 -5313 4775 -4207
rect 5423 -4340 5635 -3820
rect 6177 -3953 6239 -2847
rect 6327 -3953 6389 -2847
rect 7037 -2980 7249 -2460
rect 7791 -2593 7853 -1487
rect 7941 -2593 8003 -1487
rect 8651 -1620 8863 -1100
rect 9405 -1233 9467 -127
rect 9555 -1233 9617 -127
rect 10265 -260 10477 260
rect 11019 127 11081 1233
rect 11169 127 11231 1233
rect 11879 1100 12091 1620
rect 12633 1487 12695 2593
rect 12783 1487 12845 2593
rect 13493 2460 13705 2980
rect 14247 2847 14309 3953
rect 14397 2847 14459 3953
rect 15107 3820 15319 4340
rect 15861 4207 15923 5313
rect 16011 4207 16073 5313
rect 16721 5180 16933 5700
rect 17475 5567 17537 6673
rect 17625 5567 17687 6673
rect 17475 5313 17687 5567
rect 15861 3953 16073 4207
rect 14247 2593 14459 2847
rect 12633 1233 12845 1487
rect 11019 -127 11231 127
rect 9405 -1487 9617 -1233
rect 7791 -2847 8003 -2593
rect 6177 -4207 6389 -3953
rect 4563 -5567 4775 -5313
rect 2949 -6927 3161 -6673
rect 1335 -8160 1547 -8033
rect 2195 -8160 2407 -7900
rect 2949 -8033 3011 -6927
rect 3099 -8033 3161 -6927
rect 3809 -7060 4021 -6540
rect 4563 -6673 4625 -5567
rect 4713 -6673 4775 -5567
rect 5423 -5700 5635 -5180
rect 6177 -5313 6239 -4207
rect 6327 -5313 6389 -4207
rect 7037 -4340 7249 -3820
rect 7791 -3953 7853 -2847
rect 7941 -3953 8003 -2847
rect 8651 -2980 8863 -2460
rect 9405 -2593 9467 -1487
rect 9555 -2593 9617 -1487
rect 10265 -1620 10477 -1100
rect 11019 -1233 11081 -127
rect 11169 -1233 11231 -127
rect 11879 -260 12091 260
rect 12633 127 12695 1233
rect 12783 127 12845 1233
rect 13493 1100 13705 1620
rect 14247 1487 14309 2593
rect 14397 1487 14459 2593
rect 15107 2460 15319 2980
rect 15861 2847 15923 3953
rect 16011 2847 16073 3953
rect 16721 3820 16933 4340
rect 17475 4207 17537 5313
rect 17625 4207 17687 5313
rect 17475 3953 17687 4207
rect 15861 2593 16073 2847
rect 14247 1233 14459 1487
rect 12633 -127 12845 127
rect 11019 -1487 11231 -1233
rect 9405 -2847 9617 -2593
rect 7791 -4207 8003 -3953
rect 6177 -5567 6389 -5313
rect 4563 -6927 4775 -6673
rect 2949 -8160 3161 -8033
rect 3809 -8160 4021 -7900
rect 4563 -8033 4625 -6927
rect 4713 -8033 4775 -6927
rect 5423 -7060 5635 -6540
rect 6177 -6673 6239 -5567
rect 6327 -6673 6389 -5567
rect 7037 -5700 7249 -5180
rect 7791 -5313 7853 -4207
rect 7941 -5313 8003 -4207
rect 8651 -4340 8863 -3820
rect 9405 -3953 9467 -2847
rect 9555 -3953 9617 -2847
rect 10265 -2980 10477 -2460
rect 11019 -2593 11081 -1487
rect 11169 -2593 11231 -1487
rect 11879 -1620 12091 -1100
rect 12633 -1233 12695 -127
rect 12783 -1233 12845 -127
rect 13493 -260 13705 260
rect 14247 127 14309 1233
rect 14397 127 14459 1233
rect 15107 1100 15319 1620
rect 15861 1487 15923 2593
rect 16011 1487 16073 2593
rect 16721 2460 16933 2980
rect 17475 2847 17537 3953
rect 17625 2847 17687 3953
rect 17475 2593 17687 2847
rect 15861 1233 16073 1487
rect 14247 -127 14459 127
rect 12633 -1487 12845 -1233
rect 11019 -2847 11231 -2593
rect 9405 -4207 9617 -3953
rect 7791 -5567 8003 -5313
rect 6177 -6927 6389 -6673
rect 4563 -8160 4775 -8033
rect 5423 -8160 5635 -7900
rect 6177 -8033 6239 -6927
rect 6327 -8033 6389 -6927
rect 7037 -7060 7249 -6540
rect 7791 -6673 7853 -5567
rect 7941 -6673 8003 -5567
rect 8651 -5700 8863 -5180
rect 9405 -5313 9467 -4207
rect 9555 -5313 9617 -4207
rect 10265 -4340 10477 -3820
rect 11019 -3953 11081 -2847
rect 11169 -3953 11231 -2847
rect 11879 -2980 12091 -2460
rect 12633 -2593 12695 -1487
rect 12783 -2593 12845 -1487
rect 13493 -1620 13705 -1100
rect 14247 -1233 14309 -127
rect 14397 -1233 14459 -127
rect 15107 -260 15319 260
rect 15861 127 15923 1233
rect 16011 127 16073 1233
rect 16721 1100 16933 1620
rect 17475 1487 17537 2593
rect 17625 1487 17687 2593
rect 17475 1233 17687 1487
rect 15861 -127 16073 127
rect 14247 -1487 14459 -1233
rect 12633 -2847 12845 -2593
rect 11019 -4207 11231 -3953
rect 9405 -5567 9617 -5313
rect 7791 -6927 8003 -6673
rect 6177 -8160 6389 -8033
rect 7037 -8160 7249 -7900
rect 7791 -8033 7853 -6927
rect 7941 -8033 8003 -6927
rect 8651 -7060 8863 -6540
rect 9405 -6673 9467 -5567
rect 9555 -6673 9617 -5567
rect 10265 -5700 10477 -5180
rect 11019 -5313 11081 -4207
rect 11169 -5313 11231 -4207
rect 11879 -4340 12091 -3820
rect 12633 -3953 12695 -2847
rect 12783 -3953 12845 -2847
rect 13493 -2980 13705 -2460
rect 14247 -2593 14309 -1487
rect 14397 -2593 14459 -1487
rect 15107 -1620 15319 -1100
rect 15861 -1233 15923 -127
rect 16011 -1233 16073 -127
rect 16721 -260 16933 260
rect 17475 127 17537 1233
rect 17625 127 17687 1233
rect 17475 -127 17687 127
rect 15861 -1487 16073 -1233
rect 14247 -2847 14459 -2593
rect 12633 -4207 12845 -3953
rect 11019 -5567 11231 -5313
rect 9405 -6927 9617 -6673
rect 7791 -8160 8003 -8033
rect 8651 -8160 8863 -7900
rect 9405 -8033 9467 -6927
rect 9555 -8033 9617 -6927
rect 10265 -7060 10477 -6540
rect 11019 -6673 11081 -5567
rect 11169 -6673 11231 -5567
rect 11879 -5700 12091 -5180
rect 12633 -5313 12695 -4207
rect 12783 -5313 12845 -4207
rect 13493 -4340 13705 -3820
rect 14247 -3953 14309 -2847
rect 14397 -3953 14459 -2847
rect 15107 -2980 15319 -2460
rect 15861 -2593 15923 -1487
rect 16011 -2593 16073 -1487
rect 16721 -1620 16933 -1100
rect 17475 -1233 17537 -127
rect 17625 -1233 17687 -127
rect 17475 -1487 17687 -1233
rect 15861 -2847 16073 -2593
rect 14247 -4207 14459 -3953
rect 12633 -5567 12845 -5313
rect 11019 -6927 11231 -6673
rect 9405 -8160 9617 -8033
rect 10265 -8160 10477 -7900
rect 11019 -8033 11081 -6927
rect 11169 -8033 11231 -6927
rect 11879 -7060 12091 -6540
rect 12633 -6673 12695 -5567
rect 12783 -6673 12845 -5567
rect 13493 -5700 13705 -5180
rect 14247 -5313 14309 -4207
rect 14397 -5313 14459 -4207
rect 15107 -4340 15319 -3820
rect 15861 -3953 15923 -2847
rect 16011 -3953 16073 -2847
rect 16721 -2980 16933 -2460
rect 17475 -2593 17537 -1487
rect 17625 -2593 17687 -1487
rect 17475 -2847 17687 -2593
rect 15861 -4207 16073 -3953
rect 14247 -5567 14459 -5313
rect 12633 -6927 12845 -6673
rect 11019 -8160 11231 -8033
rect 11879 -8160 12091 -7900
rect 12633 -8033 12695 -6927
rect 12783 -8033 12845 -6927
rect 13493 -7060 13705 -6540
rect 14247 -6673 14309 -5567
rect 14397 -6673 14459 -5567
rect 15107 -5700 15319 -5180
rect 15861 -5313 15923 -4207
rect 16011 -5313 16073 -4207
rect 16721 -4340 16933 -3820
rect 17475 -3953 17537 -2847
rect 17625 -3953 17687 -2847
rect 17475 -4207 17687 -3953
rect 15861 -5567 16073 -5313
rect 14247 -6927 14459 -6673
rect 12633 -8160 12845 -8033
rect 13493 -8160 13705 -7900
rect 14247 -8033 14309 -6927
rect 14397 -8033 14459 -6927
rect 15107 -7060 15319 -6540
rect 15861 -6673 15923 -5567
rect 16011 -6673 16073 -5567
rect 16721 -5700 16933 -5180
rect 17475 -5313 17537 -4207
rect 17625 -5313 17687 -4207
rect 17475 -5567 17687 -5313
rect 15861 -6927 16073 -6673
rect 14247 -8160 14459 -8033
rect 15107 -8160 15319 -7900
rect 15861 -8033 15923 -6927
rect 16011 -8033 16073 -6927
rect 16721 -7060 16933 -6540
rect 17475 -6673 17537 -5567
rect 17625 -6673 17687 -5567
rect 17475 -6927 17687 -6673
rect 15861 -8160 16073 -8033
rect 16721 -8160 16933 -7900
rect 17475 -8033 17537 -6927
rect 17625 -8033 17687 -6927
rect 17475 -8160 17687 -8033
<< properties >>
string FIXED_BBOX 16207 6860 17447 8100
string gencell cap_mim_2p0fF
string library gf180mcu
string parameters w 5.00 l 5.00 val 1.025k carea 25.00 cperi 20.00 class capacitor nx 22 ny 12 dummy 0 square 0 lmin 5.00 wmin 5.00 lmax 100.0 wmax 100.0 dc 0 bconnect 1 tconnect 1
<< end >>
