magic
tech gf180mcuD
magscale 1 10
timestamp 1755276408
<< pwell >>
rect -336 -15456 336 15456
<< psubdiff >>
rect -312 15360 312 15432
rect -312 15316 -240 15360
rect -312 -15316 -299 15316
rect -253 -15316 -240 15316
rect 240 15316 312 15360
rect -312 -15360 -240 -15316
rect 240 -15316 253 15316
rect 299 -15316 312 15316
rect 240 -15360 312 -15316
rect -312 -15432 312 -15360
<< psubdiffcont >>
rect -299 -15316 -253 15316
rect 253 -15316 299 15316
<< polysilicon >>
rect -100 15207 100 15220
rect -100 15161 -87 15207
rect 87 15161 100 15207
rect -100 15098 100 15161
rect -100 12361 100 12424
rect -100 12315 -87 12361
rect 87 12315 100 12361
rect -100 12302 100 12315
rect -100 12149 100 12162
rect -100 12103 -87 12149
rect 87 12103 100 12149
rect -100 12040 100 12103
rect -100 9303 100 9366
rect -100 9257 -87 9303
rect 87 9257 100 9303
rect -100 9244 100 9257
rect -100 9091 100 9104
rect -100 9045 -87 9091
rect 87 9045 100 9091
rect -100 8982 100 9045
rect -100 6245 100 6308
rect -100 6199 -87 6245
rect 87 6199 100 6245
rect -100 6186 100 6199
rect -100 6033 100 6046
rect -100 5987 -87 6033
rect 87 5987 100 6033
rect -100 5924 100 5987
rect -100 3187 100 3250
rect -100 3141 -87 3187
rect 87 3141 100 3187
rect -100 3128 100 3141
rect -100 2975 100 2988
rect -100 2929 -87 2975
rect 87 2929 100 2975
rect -100 2866 100 2929
rect -100 129 100 192
rect -100 83 -87 129
rect 87 83 100 129
rect -100 70 100 83
rect -100 -83 100 -70
rect -100 -129 -87 -83
rect 87 -129 100 -83
rect -100 -192 100 -129
rect -100 -2929 100 -2866
rect -100 -2975 -87 -2929
rect 87 -2975 100 -2929
rect -100 -2988 100 -2975
rect -100 -3141 100 -3128
rect -100 -3187 -87 -3141
rect 87 -3187 100 -3141
rect -100 -3250 100 -3187
rect -100 -5987 100 -5924
rect -100 -6033 -87 -5987
rect 87 -6033 100 -5987
rect -100 -6046 100 -6033
rect -100 -6199 100 -6186
rect -100 -6245 -87 -6199
rect 87 -6245 100 -6199
rect -100 -6308 100 -6245
rect -100 -9045 100 -8982
rect -100 -9091 -87 -9045
rect 87 -9091 100 -9045
rect -100 -9104 100 -9091
rect -100 -9257 100 -9244
rect -100 -9303 -87 -9257
rect 87 -9303 100 -9257
rect -100 -9366 100 -9303
rect -100 -12103 100 -12040
rect -100 -12149 -87 -12103
rect 87 -12149 100 -12103
rect -100 -12162 100 -12149
rect -100 -12315 100 -12302
rect -100 -12361 -87 -12315
rect 87 -12361 100 -12315
rect -100 -12424 100 -12361
rect -100 -15161 100 -15098
rect -100 -15207 -87 -15161
rect 87 -15207 100 -15161
rect -100 -15220 100 -15207
<< polycontact >>
rect -87 15161 87 15207
rect -87 12315 87 12361
rect -87 12103 87 12149
rect -87 9257 87 9303
rect -87 9045 87 9091
rect -87 6199 87 6245
rect -87 5987 87 6033
rect -87 3141 87 3187
rect -87 2929 87 2975
rect -87 83 87 129
rect -87 -129 87 -83
rect -87 -2975 87 -2929
rect -87 -3187 87 -3141
rect -87 -6033 87 -5987
rect -87 -6245 87 -6199
rect -87 -9091 87 -9045
rect -87 -9303 87 -9257
rect -87 -12149 87 -12103
rect -87 -12361 87 -12315
rect -87 -15207 87 -15161
<< nhighres >>
rect -100 12424 100 15098
rect -100 9366 100 12040
rect -100 6308 100 8982
rect -100 3250 100 5924
rect -100 192 100 2866
rect -100 -2866 100 -192
rect -100 -5924 100 -3250
rect -100 -8982 100 -6308
rect -100 -12040 100 -9366
rect -100 -15098 100 -12424
<< metal1 >>
rect -299 15373 299 15419
rect -299 15316 -253 15373
rect 253 15316 299 15373
rect -98 15161 -87 15207
rect 87 15161 98 15207
rect -98 12315 -87 12361
rect 87 12315 98 12361
rect -98 12103 -87 12149
rect 87 12103 98 12149
rect -98 9257 -87 9303
rect 87 9257 98 9303
rect -98 9045 -87 9091
rect 87 9045 98 9091
rect -98 6199 -87 6245
rect 87 6199 98 6245
rect -98 5987 -87 6033
rect 87 5987 98 6033
rect -98 3141 -87 3187
rect 87 3141 98 3187
rect -98 2929 -87 2975
rect 87 2929 98 2975
rect -98 83 -87 129
rect 87 83 98 129
rect -98 -129 -87 -83
rect 87 -129 98 -83
rect -98 -2975 -87 -2929
rect 87 -2975 98 -2929
rect -98 -3187 -87 -3141
rect 87 -3187 98 -3141
rect -98 -6033 -87 -5987
rect 87 -6033 98 -5987
rect -98 -6245 -87 -6199
rect 87 -6245 98 -6199
rect -98 -9091 -87 -9045
rect 87 -9091 98 -9045
rect -98 -9303 -87 -9257
rect 87 -9303 98 -9257
rect -98 -12149 -87 -12103
rect 87 -12149 98 -12103
rect -98 -12361 -87 -12315
rect 87 -12361 98 -12315
rect -98 -15207 -87 -15161
rect 87 -15207 98 -15161
rect -299 -15373 -253 -15316
rect 253 -15373 299 -15316
rect -299 -15419 299 -15373
<< properties >>
string FIXED_BBOX -276 -15396 276 15396
string gencell ppolyf_u_1k
string library gf180mcu
string parameters w 1.0 l 13.37 m 10 nx 1 wmin 1.000 lmin 1.000 class resistor rho 1000 val 13.37k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
