magic
tech gf180mcuD
magscale 1 5
timestamp 1757579644
<< checkpaint >>
rect -1030 -1430 1286 988
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
use ppolyf_u_EJ86NH  XR1
timestamp 0
transform 1 0 128 0 1 -221
box -158 -209 158 209
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 640 0 0 0 A
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 640 0 0 0 B
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 640 0 0 0 C
port 2 nsew
<< end >>
